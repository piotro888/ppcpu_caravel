magic
tech sky130B
magscale 1 2
timestamp 1663051890
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 235166 700612 235172 700664
rect 235224 700652 235230 700664
rect 253290 700652 253296 700664
rect 235224 700624 253296 700652
rect 235224 700612 235230 700624
rect 253290 700612 253296 700624
rect 253348 700612 253354 700664
rect 218974 700544 218980 700596
rect 219032 700584 219038 700596
rect 253382 700584 253388 700596
rect 219032 700556 253388 700584
rect 219032 700544 219038 700556
rect 253382 700544 253388 700556
rect 253440 700544 253446 700596
rect 154114 700476 154120 700528
rect 154172 700516 154178 700528
rect 264330 700516 264336 700528
rect 154172 700488 264336 700516
rect 154172 700476 154178 700488
rect 264330 700476 264336 700488
rect 264388 700476 264394 700528
rect 283834 700476 283840 700528
rect 283892 700516 283898 700528
rect 477034 700516 477040 700528
rect 283892 700488 477040 700516
rect 283892 700476 283898 700488
rect 477034 700476 477040 700488
rect 477092 700476 477098 700528
rect 89162 700408 89168 700460
rect 89220 700448 89226 700460
rect 265618 700448 265624 700460
rect 89220 700420 265624 700448
rect 89220 700408 89226 700420
rect 265618 700408 265624 700420
rect 265676 700408 265682 700460
rect 300118 700408 300124 700460
rect 300176 700448 300182 700460
rect 320910 700448 320916 700460
rect 300176 700420 320916 700448
rect 300176 700408 300182 700420
rect 320910 700408 320916 700420
rect 320968 700408 320974 700460
rect 360838 700408 360844 700460
rect 360896 700448 360902 700460
rect 559650 700448 559656 700460
rect 360896 700420 559656 700448
rect 360896 700408 360902 700420
rect 559650 700408 559656 700420
rect 559708 700408 559714 700460
rect 72970 700340 72976 700392
rect 73028 700380 73034 700392
rect 253198 700380 253204 700392
rect 73028 700352 253204 700380
rect 73028 700340 73034 700352
rect 253198 700340 253204 700352
rect 253256 700340 253262 700392
rect 317414 700340 317420 700392
rect 317472 700380 317478 700392
rect 543458 700380 543464 700392
rect 317472 700352 543464 700380
rect 317472 700340 317478 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 406378 700312 406384 700324
rect 24360 700284 406384 700312
rect 24360 700272 24366 700284
rect 406378 700272 406384 700284
rect 406436 700272 406442 700324
rect 520918 699660 520924 699712
rect 520976 699700 520982 699712
rect 527174 699700 527180 699712
rect 520976 699672 527180 699700
rect 520976 699660 520982 699672
rect 527174 699660 527180 699672
rect 527232 699660 527238 699712
rect 397454 698912 397460 698964
rect 397512 698952 397518 698964
rect 477126 698952 477132 698964
rect 397512 698924 477132 698952
rect 397512 698912 397518 698924
rect 477126 698912 477132 698924
rect 477184 698912 477190 698964
rect 266354 697620 266360 697672
rect 266412 697660 266418 697672
rect 267642 697660 267648 697672
rect 266412 697632 267648 697660
rect 266412 697620 266418 697632
rect 267642 697620 267648 697632
rect 267700 697620 267706 697672
rect 105446 697552 105452 697604
rect 105504 697592 105510 697604
rect 337378 697592 337384 697604
rect 105504 697564 337384 697592
rect 105504 697552 105510 697564
rect 337378 697552 337384 697564
rect 337436 697552 337442 697604
rect 525150 696940 525156 696992
rect 525208 696980 525214 696992
rect 580166 696980 580172 696992
rect 525208 696952 580172 696980
rect 525208 696940 525214 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 316126 683136 316132 683188
rect 316184 683176 316190 683188
rect 580166 683176 580172 683188
rect 316184 683148 580172 683176
rect 316184 683136 316190 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 403710 670692 403716 670744
rect 403768 670732 403774 670744
rect 580166 670732 580172 670744
rect 403768 670704 580172 670732
rect 403768 670692 403774 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 6914 665796 6920 665848
rect 6972 665836 6978 665848
rect 475746 665836 475752 665848
rect 6972 665808 475752 665836
rect 6972 665796 6978 665808
rect 475746 665796 475752 665808
rect 475804 665796 475810 665848
rect 52086 663824 52092 663876
rect 52144 663864 52150 663876
rect 355410 663864 355416 663876
rect 52144 663836 355416 663864
rect 52144 663824 52150 663836
rect 355410 663824 355416 663836
rect 355468 663824 355474 663876
rect 46474 663756 46480 663808
rect 46532 663796 46538 663808
rect 352558 663796 352564 663808
rect 46532 663768 352564 663796
rect 46532 663756 46538 663768
rect 352558 663756 352564 663768
rect 352616 663756 352622 663808
rect 50430 663076 50436 663128
rect 50488 663116 50494 663128
rect 279418 663116 279424 663128
rect 50488 663088 279424 663116
rect 50488 663076 50494 663088
rect 279418 663076 279424 663088
rect 279476 663076 279482 663128
rect 46750 663008 46756 663060
rect 46808 663048 46814 663060
rect 279970 663048 279976 663060
rect 46808 663020 279976 663048
rect 46808 663008 46814 663020
rect 279970 663008 279976 663020
rect 280028 663008 280034 663060
rect 51718 662940 51724 662992
rect 51776 662980 51782 662992
rect 352834 662980 352840 662992
rect 51776 662952 352840 662980
rect 51776 662940 51782 662952
rect 352834 662940 352840 662952
rect 352892 662940 352898 662992
rect 51074 662872 51080 662924
rect 51132 662912 51138 662924
rect 352650 662912 352656 662924
rect 51132 662884 352656 662912
rect 51132 662872 51138 662884
rect 352650 662872 352656 662884
rect 352708 662872 352714 662924
rect 50890 662804 50896 662856
rect 50948 662844 50954 662856
rect 353018 662844 353024 662856
rect 50948 662816 353024 662844
rect 50948 662804 50954 662816
rect 353018 662804 353024 662816
rect 353076 662804 353082 662856
rect 51994 662736 52000 662788
rect 52052 662776 52058 662788
rect 355318 662776 355324 662788
rect 52052 662748 355324 662776
rect 52052 662736 52058 662748
rect 355318 662736 355324 662748
rect 355376 662736 355382 662788
rect 47854 662668 47860 662720
rect 47912 662708 47918 662720
rect 352926 662708 352932 662720
rect 47912 662680 352932 662708
rect 47912 662668 47918 662680
rect 352926 662668 352932 662680
rect 352984 662668 352990 662720
rect 45462 662600 45468 662652
rect 45520 662640 45526 662652
rect 352742 662640 352748 662652
rect 45520 662612 352748 662640
rect 45520 662600 45526 662612
rect 352742 662600 352748 662612
rect 352800 662600 352806 662652
rect 51902 662532 51908 662584
rect 51960 662572 51966 662584
rect 405090 662572 405096 662584
rect 51960 662544 405096 662572
rect 51960 662532 51966 662544
rect 405090 662532 405096 662544
rect 405148 662532 405154 662584
rect 52178 662464 52184 662516
rect 52236 662504 52242 662516
rect 405734 662504 405740 662516
rect 52236 662476 405740 662504
rect 52236 662464 52242 662476
rect 405734 662464 405740 662476
rect 405792 662464 405798 662516
rect 46382 662396 46388 662448
rect 46440 662436 46446 662448
rect 403802 662436 403808 662448
rect 46440 662408 403808 662436
rect 46440 662396 46446 662408
rect 403802 662396 403808 662408
rect 403860 662396 403866 662448
rect 201494 661784 201500 661836
rect 201552 661824 201558 661836
rect 422938 661824 422944 661836
rect 201552 661796 422944 661824
rect 201552 661784 201558 661796
rect 422938 661784 422944 661796
rect 422996 661784 423002 661836
rect 50246 661716 50252 661768
rect 50304 661756 50310 661768
rect 279326 661756 279332 661768
rect 50304 661728 279332 661756
rect 50304 661716 50310 661728
rect 279326 661716 279332 661728
rect 279384 661716 279390 661768
rect 136634 661648 136640 661700
rect 136692 661688 136698 661700
rect 475654 661688 475660 661700
rect 136692 661660 475660 661688
rect 136692 661648 136698 661660
rect 475654 661648 475660 661660
rect 475712 661648 475718 661700
rect 50522 661580 50528 661632
rect 50580 661620 50586 661632
rect 280062 661620 280068 661632
rect 50580 661592 280068 661620
rect 50580 661580 50586 661592
rect 280062 661580 280068 661592
rect 280120 661580 280126 661632
rect 49142 661512 49148 661564
rect 49200 661552 49206 661564
rect 279510 661552 279516 661564
rect 49200 661524 279516 661552
rect 49200 661512 49206 661524
rect 279510 661512 279516 661524
rect 279568 661512 279574 661564
rect 50798 661444 50804 661496
rect 50856 661484 50862 661496
rect 356882 661484 356888 661496
rect 50856 661456 356888 661484
rect 50856 661444 50862 661456
rect 356882 661444 356888 661456
rect 356940 661444 356946 661496
rect 50614 661376 50620 661428
rect 50672 661416 50678 661428
rect 401594 661416 401600 661428
rect 50672 661388 401600 661416
rect 50672 661376 50678 661388
rect 401594 661376 401600 661388
rect 401652 661376 401658 661428
rect 51810 661308 51816 661360
rect 51868 661348 51874 661360
rect 405826 661348 405832 661360
rect 51868 661320 405832 661348
rect 51868 661308 51874 661320
rect 405826 661308 405832 661320
rect 405884 661308 405890 661360
rect 49786 661240 49792 661292
rect 49844 661280 49850 661292
rect 511994 661280 512000 661292
rect 49844 661252 512000 661280
rect 49844 661240 49850 661252
rect 511994 661240 512000 661252
rect 512052 661240 512058 661292
rect 3602 661172 3608 661224
rect 3660 661212 3666 661224
rect 478874 661212 478880 661224
rect 3660 661184 478880 661212
rect 3660 661172 3666 661184
rect 478874 661172 478880 661184
rect 478932 661172 478938 661224
rect 3418 661104 3424 661156
rect 3476 661144 3482 661156
rect 484394 661144 484400 661156
rect 3476 661116 484400 661144
rect 3476 661104 3482 661116
rect 484394 661104 484400 661116
rect 484452 661104 484458 661156
rect 3786 661036 3792 661088
rect 3844 661076 3850 661088
rect 498194 661076 498200 661088
rect 3844 661048 498200 661076
rect 3844 661036 3850 661048
rect 498194 661036 498200 661048
rect 498252 661036 498258 661088
rect 49418 660560 49424 660612
rect 49476 660600 49482 660612
rect 257430 660600 257436 660612
rect 49476 660572 257436 660600
rect 49476 660560 49482 660572
rect 257430 660560 257436 660572
rect 257488 660560 257494 660612
rect 49602 660492 49608 660544
rect 49660 660532 49666 660544
rect 278130 660532 278136 660544
rect 49660 660504 278136 660532
rect 49660 660492 49666 660504
rect 278130 660492 278136 660504
rect 278188 660492 278194 660544
rect 50154 660424 50160 660476
rect 50212 660464 50218 660476
rect 488534 660464 488540 660476
rect 50212 660436 488540 660464
rect 50212 660424 50218 660436
rect 488534 660424 488540 660436
rect 488592 660424 488598 660476
rect 50706 660356 50712 660408
rect 50764 660396 50770 660408
rect 279602 660396 279608 660408
rect 50764 660368 279608 660396
rect 50764 660356 50770 660368
rect 279602 660356 279608 660368
rect 279660 660356 279666 660408
rect 50338 660288 50344 660340
rect 50396 660328 50402 660340
rect 500954 660328 500960 660340
rect 50396 660300 500960 660328
rect 50396 660288 50402 660300
rect 500954 660288 500960 660300
rect 501012 660288 501018 660340
rect 49510 660220 49516 660272
rect 49568 660260 49574 660272
rect 279050 660260 279056 660272
rect 49568 660232 279056 660260
rect 49568 660220 49574 660232
rect 279050 660220 279056 660232
rect 279108 660220 279114 660272
rect 49234 660152 49240 660204
rect 49292 660192 49298 660204
rect 279142 660192 279148 660204
rect 49292 660164 279148 660192
rect 49292 660152 49298 660164
rect 279142 660152 279148 660164
rect 279200 660152 279206 660204
rect 48222 660084 48228 660136
rect 48280 660124 48286 660136
rect 278958 660124 278964 660136
rect 48280 660096 278964 660124
rect 48280 660084 48286 660096
rect 278958 660084 278964 660096
rect 279016 660084 279022 660136
rect 46842 660016 46848 660068
rect 46900 660056 46906 660068
rect 279234 660056 279240 660068
rect 46900 660028 279240 660056
rect 46900 660016 46906 660028
rect 279234 660016 279240 660028
rect 279292 660016 279298 660068
rect 51350 659948 51356 660000
rect 51408 659988 51414 660000
rect 296898 659988 296904 660000
rect 51408 659960 296904 659988
rect 51408 659948 51414 659960
rect 296898 659948 296904 659960
rect 296956 659948 296962 660000
rect 51258 659880 51264 659932
rect 51316 659920 51322 659932
rect 356974 659920 356980 659932
rect 51316 659892 356980 659920
rect 51316 659880 51322 659892
rect 356974 659880 356980 659892
rect 357032 659880 357038 659932
rect 3326 659812 3332 659864
rect 3384 659852 3390 659864
rect 477218 659852 477224 659864
rect 3384 659824 477224 659852
rect 3384 659812 3390 659824
rect 477218 659812 477224 659824
rect 477276 659812 477282 659864
rect 50338 658656 50344 658708
rect 50396 658696 50402 658708
rect 50982 658696 50988 658708
rect 50396 658668 50988 658696
rect 50396 658656 50402 658668
rect 50982 658656 50988 658668
rect 51040 658656 51046 658708
rect 254578 656888 254584 656940
rect 254636 656928 254642 656940
rect 353110 656928 353116 656940
rect 254636 656900 353116 656928
rect 254636 656888 254642 656900
rect 353110 656888 353116 656900
rect 353168 656888 353174 656940
rect 48682 652740 48688 652792
rect 48740 652780 48746 652792
rect 49970 652780 49976 652792
rect 48740 652752 49976 652780
rect 48740 652740 48746 652752
rect 49970 652740 49976 652752
rect 50028 652740 50034 652792
rect 50982 651380 50988 651432
rect 51040 651420 51046 651432
rect 52178 651420 52184 651432
rect 51040 651392 52184 651420
rect 51040 651380 51046 651392
rect 52178 651380 52184 651392
rect 52236 651380 52242 651432
rect 49234 648524 49240 648576
rect 49292 648564 49298 648576
rect 50154 648564 50160 648576
rect 49292 648536 50160 648564
rect 49292 648524 49298 648536
rect 50154 648524 50160 648536
rect 50212 648524 50218 648576
rect 253934 645872 253940 645924
rect 253992 645912 253998 645924
rect 257338 645912 257344 645924
rect 253992 645884 257344 645912
rect 253992 645872 253998 645884
rect 257338 645872 257344 645884
rect 257396 645872 257402 645924
rect 526438 643084 526444 643136
rect 526496 643124 526502 643136
rect 580166 643124 580172 643136
rect 526496 643096 580172 643124
rect 526496 643084 526502 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 357342 642812 357348 642864
rect 357400 642852 357406 642864
rect 371694 642852 371700 642864
rect 357400 642824 371700 642852
rect 357400 642812 357406 642824
rect 371694 642812 371700 642824
rect 371752 642812 371758 642864
rect 361022 642744 361028 642796
rect 361080 642784 361086 642796
rect 379974 642784 379980 642796
rect 361080 642756 379980 642784
rect 361080 642744 361086 642756
rect 379974 642744 379980 642756
rect 380032 642744 380038 642796
rect 353202 642676 353208 642728
rect 353260 642716 353266 642728
rect 382182 642716 382188 642728
rect 353260 642688 382188 642716
rect 353260 642676 353266 642688
rect 382182 642676 382188 642688
rect 382240 642676 382246 642728
rect 357250 642608 357256 642660
rect 357308 642648 357314 642660
rect 388806 642648 388812 642660
rect 357308 642620 388812 642648
rect 357308 642608 357314 642620
rect 388806 642608 388812 642620
rect 388864 642608 388870 642660
rect 392670 642608 392676 642660
rect 392728 642648 392734 642660
rect 399294 642648 399300 642660
rect 392728 642620 399300 642648
rect 392728 642608 392734 642620
rect 399294 642608 399300 642620
rect 399352 642608 399358 642660
rect 359458 642540 359464 642592
rect 359516 642580 359522 642592
rect 376110 642580 376116 642592
rect 359516 642552 376116 642580
rect 359516 642540 359522 642552
rect 376110 642540 376116 642552
rect 376168 642540 376174 642592
rect 376202 642540 376208 642592
rect 376260 642580 376266 642592
rect 400306 642580 400312 642592
rect 376260 642552 400312 642580
rect 376260 642540 376266 642552
rect 400306 642540 400312 642552
rect 400364 642540 400370 642592
rect 370038 642472 370044 642524
rect 370096 642512 370102 642524
rect 403158 642512 403164 642524
rect 370096 642484 403164 642512
rect 370096 642472 370102 642484
rect 403158 642472 403164 642484
rect 403216 642472 403222 642524
rect 310422 642404 310428 642456
rect 310480 642444 310486 642456
rect 361758 642444 361764 642456
rect 310480 642416 361764 642444
rect 310480 642404 310486 642416
rect 361758 642404 361764 642416
rect 361816 642404 361822 642456
rect 366174 642404 366180 642456
rect 366232 642444 366238 642456
rect 399110 642444 399116 642456
rect 366232 642416 399116 642444
rect 366232 642404 366238 642416
rect 399110 642404 399116 642416
rect 399168 642404 399174 642456
rect 287606 642336 287612 642388
rect 287664 642376 287670 642388
rect 351362 642376 351368 642388
rect 287664 642348 351368 642376
rect 287664 642336 287670 642348
rect 351362 642336 351368 642348
rect 351420 642336 351426 642388
rect 355962 642336 355968 642388
rect 356020 642376 356026 642388
rect 391014 642376 391020 642388
rect 356020 642348 391020 642376
rect 356020 642336 356026 642348
rect 391014 642336 391020 642348
rect 391072 642336 391078 642388
rect 392118 642336 392124 642388
rect 392176 642376 392182 642388
rect 399202 642376 399208 642388
rect 392176 642348 399208 642376
rect 392176 642336 392182 642348
rect 399202 642336 399208 642348
rect 399260 642336 399266 642388
rect 293126 642268 293132 642320
rect 293184 642308 293190 642320
rect 321094 642308 321100 642320
rect 293184 642280 321100 642308
rect 293184 642268 293190 642280
rect 321094 642268 321100 642280
rect 321152 642268 321158 642320
rect 365530 642268 365536 642320
rect 365588 642308 365594 642320
rect 383286 642308 383292 642320
rect 365588 642280 383292 642308
rect 365588 642268 365594 642280
rect 383286 642268 383292 642280
rect 383344 642268 383350 642320
rect 393222 642268 393228 642320
rect 393280 642308 393286 642320
rect 400490 642308 400496 642320
rect 393280 642280 400496 642308
rect 393280 642268 393286 642280
rect 400490 642268 400496 642280
rect 400548 642268 400554 642320
rect 295242 642200 295248 642252
rect 295300 642240 295306 642252
rect 323670 642240 323676 642252
rect 295300 642212 323676 642240
rect 295300 642200 295306 642212
rect 323670 642200 323676 642212
rect 323728 642200 323734 642252
rect 349890 642200 349896 642252
rect 349948 642240 349954 642252
rect 377766 642240 377772 642252
rect 349948 642212 377772 642240
rect 349948 642200 349954 642212
rect 377766 642200 377772 642212
rect 377824 642200 377830 642252
rect 387150 642200 387156 642252
rect 387208 642240 387214 642252
rect 400950 642240 400956 642252
rect 387208 642212 400956 642240
rect 387208 642200 387214 642212
rect 400950 642200 400956 642212
rect 401008 642200 401014 642252
rect 300762 642132 300768 642184
rect 300820 642172 300826 642184
rect 329190 642172 329196 642184
rect 300820 642144 329196 642172
rect 300820 642132 300826 642144
rect 329190 642132 329196 642144
rect 329248 642132 329254 642184
rect 355594 642132 355600 642184
rect 355652 642172 355658 642184
rect 386046 642172 386052 642184
rect 355652 642144 386052 642172
rect 355652 642132 355658 642144
rect 386046 642132 386052 642144
rect 386104 642132 386110 642184
rect 394326 642132 394332 642184
rect 394384 642172 394390 642184
rect 405274 642172 405280 642184
rect 394384 642144 405280 642172
rect 394384 642132 394390 642144
rect 405274 642132 405280 642144
rect 405332 642132 405338 642184
rect 286502 642064 286508 642116
rect 286560 642104 286566 642116
rect 321002 642104 321008 642116
rect 286560 642076 321008 642104
rect 286560 642064 286566 642076
rect 321002 642064 321008 642076
rect 321060 642064 321066 642116
rect 371142 642064 371148 642116
rect 371200 642104 371206 642116
rect 399662 642104 399668 642116
rect 371200 642076 399668 642104
rect 371200 642064 371206 642076
rect 399662 642064 399668 642076
rect 399720 642064 399726 642116
rect 296346 641996 296352 642048
rect 296404 642036 296410 642048
rect 331858 642036 331864 642048
rect 296404 642008 331864 642036
rect 296404 641996 296410 642008
rect 331858 641996 331864 642008
rect 331916 641996 331922 642048
rect 333238 641996 333244 642048
rect 333296 642036 333302 642048
rect 363414 642036 363420 642048
rect 333296 642008 363420 642036
rect 333296 641996 333302 642008
rect 363414 641996 363420 642008
rect 363472 641996 363478 642048
rect 374454 641996 374460 642048
rect 374512 642036 374518 642048
rect 405182 642036 405188 642048
rect 374512 642008 405188 642036
rect 374512 641996 374518 642008
rect 405182 641996 405188 642008
rect 405240 641996 405246 642048
rect 284202 641928 284208 641980
rect 284260 641968 284266 641980
rect 325050 641968 325056 641980
rect 284260 641940 325056 641968
rect 284260 641928 284266 641940
rect 325050 641928 325056 641940
rect 325108 641928 325114 641980
rect 359734 641928 359740 641980
rect 359792 641968 359798 641980
rect 373350 641968 373356 641980
rect 359792 641940 373356 641968
rect 359792 641928 359798 641940
rect 373350 641928 373356 641940
rect 373408 641928 373414 641980
rect 290918 641860 290924 641912
rect 290976 641900 290982 641912
rect 319438 641900 319444 641912
rect 290976 641872 319444 641900
rect 290976 641860 290982 641872
rect 319438 641860 319444 641872
rect 319496 641860 319502 641912
rect 357066 641860 357072 641912
rect 357124 641900 357130 641912
rect 381078 641900 381084 641912
rect 357124 641872 381084 641900
rect 357124 641860 357130 641872
rect 381078 641860 381084 641872
rect 381136 641860 381142 641912
rect 394878 641860 394884 641912
rect 394936 641900 394942 641912
rect 400582 641900 400588 641912
rect 394936 641872 400588 641900
rect 394936 641860 394942 641872
rect 400582 641860 400588 641872
rect 400640 641860 400646 641912
rect 297542 641792 297548 641844
rect 297600 641832 297606 641844
rect 349798 641832 349804 641844
rect 297600 641804 349804 641832
rect 297600 641792 297606 641804
rect 349798 641792 349804 641804
rect 349856 641792 349862 641844
rect 360102 641792 360108 641844
rect 360160 641832 360166 641844
rect 368382 641832 368388 641844
rect 360160 641804 368388 641832
rect 360160 641792 360166 641804
rect 368382 641792 368388 641804
rect 368440 641792 368446 641844
rect 378042 641792 378048 641844
rect 378100 641832 378106 641844
rect 386598 641832 386604 641844
rect 378100 641804 386604 641832
rect 378100 641792 378106 641804
rect 386598 641792 386604 641804
rect 386656 641792 386662 641844
rect 393774 641792 393780 641844
rect 393832 641832 393838 641844
rect 399386 641832 399392 641844
rect 393832 641804 399392 641832
rect 393832 641792 393838 641804
rect 399386 641792 399392 641804
rect 399444 641792 399450 641844
rect 472618 641792 472624 641844
rect 472676 641832 472682 641844
rect 493226 641832 493232 641844
rect 472676 641804 493232 641832
rect 472676 641792 472682 641804
rect 493226 641792 493232 641804
rect 493284 641792 493290 641844
rect 49050 641724 49056 641776
rect 49108 641764 49114 641776
rect 50246 641764 50252 641776
rect 49108 641736 50252 641764
rect 49108 641724 49114 641736
rect 50246 641724 50252 641736
rect 50304 641724 50310 641776
rect 358814 641724 358820 641776
rect 358872 641764 358878 641776
rect 366726 641764 366732 641776
rect 358872 641736 366732 641764
rect 358872 641724 358878 641736
rect 366726 641724 366732 641736
rect 366784 641724 366790 641776
rect 375558 641724 375564 641776
rect 375616 641764 375622 641776
rect 376202 641764 376208 641776
rect 375616 641736 376208 641764
rect 375616 641724 375622 641736
rect 376202 641724 376208 641736
rect 376260 641724 376266 641776
rect 395430 641724 395436 641776
rect 395488 641764 395494 641776
rect 399754 641764 399760 641776
rect 395488 641736 399760 641764
rect 395488 641724 395494 641736
rect 399754 641724 399760 641736
rect 399812 641724 399818 641776
rect 404998 641724 405004 641776
rect 405056 641764 405062 641776
rect 510614 641764 510620 641776
rect 405056 641736 510620 641764
rect 405056 641724 405062 641736
rect 510614 641724 510620 641736
rect 510672 641724 510678 641776
rect 358538 641180 358544 641232
rect 358596 641220 358602 641232
rect 391566 641220 391572 641232
rect 358596 641192 391572 641220
rect 358596 641180 358602 641192
rect 391566 641180 391572 641192
rect 391624 641180 391630 641232
rect 278682 641112 278688 641164
rect 278740 641152 278746 641164
rect 398466 641152 398472 641164
rect 278740 641124 398472 641152
rect 278740 641112 278746 641124
rect 398466 641112 398472 641124
rect 398524 641112 398530 641164
rect 315850 641044 315856 641096
rect 315908 641084 315914 641096
rect 523678 641084 523684 641096
rect 315908 641056 523684 641084
rect 315908 641044 315914 641056
rect 523678 641044 523684 641056
rect 523736 641044 523742 641096
rect 278590 640976 278596 641028
rect 278648 641016 278654 641028
rect 310422 641016 310428 641028
rect 278648 640988 310428 641016
rect 278648 640976 278654 640988
rect 310422 640976 310428 640988
rect 310480 640976 310486 641028
rect 314102 640976 314108 641028
rect 314160 641016 314166 641028
rect 530578 641016 530584 641028
rect 314160 640988 530584 641016
rect 314160 640976 314166 640988
rect 530578 640976 530584 640988
rect 530636 640976 530642 641028
rect 355502 640908 355508 640960
rect 355560 640948 355566 640960
rect 378318 640948 378324 640960
rect 355560 640920 378324 640948
rect 355560 640908 355566 640920
rect 378318 640908 378324 640920
rect 378376 640908 378382 640960
rect 357158 640840 357164 640892
rect 357216 640880 357222 640892
rect 383838 640880 383844 640892
rect 357216 640852 383844 640880
rect 357216 640840 357222 640852
rect 383838 640840 383844 640852
rect 383896 640840 383902 640892
rect 357802 640772 357808 640824
rect 357860 640812 357866 640824
rect 388254 640812 388260 640824
rect 357860 640784 388260 640812
rect 357860 640772 357866 640784
rect 388254 640772 388260 640784
rect 388312 640772 388318 640824
rect 359182 640704 359188 640756
rect 359240 640744 359246 640756
rect 389358 640744 389364 640756
rect 359240 640716 389364 640744
rect 359240 640704 359246 640716
rect 389358 640704 389364 640716
rect 389416 640704 389422 640756
rect 312998 640636 313004 640688
rect 313056 640676 313062 640688
rect 338758 640676 338764 640688
rect 313056 640648 338764 640676
rect 313056 640636 313062 640648
rect 338758 640636 338764 640648
rect 338816 640636 338822 640688
rect 342898 640636 342904 640688
rect 342956 640676 342962 640688
rect 384942 640676 384948 640688
rect 342956 640648 384948 640676
rect 342956 640636 342962 640648
rect 384942 640636 384948 640648
rect 385000 640636 385006 640688
rect 387702 640636 387708 640688
rect 387760 640676 387766 640688
rect 401870 640676 401876 640688
rect 387760 640648 401876 640676
rect 387760 640636 387766 640648
rect 401870 640636 401876 640648
rect 401928 640636 401934 640688
rect 308582 640568 308588 640620
rect 308640 640608 308646 640620
rect 356790 640608 356796 640620
rect 308640 640580 356796 640608
rect 308640 640568 308646 640580
rect 356790 640568 356796 640580
rect 356848 640568 356854 640620
rect 389910 640568 389916 640620
rect 389968 640608 389974 640620
rect 401594 640608 401600 640620
rect 389968 640580 401600 640608
rect 389968 640568 389974 640580
rect 401594 640568 401600 640580
rect 401652 640568 401658 640620
rect 303062 640500 303068 640552
rect 303120 640540 303126 640552
rect 356698 640540 356704 640552
rect 303120 640512 356704 640540
rect 303120 640500 303126 640512
rect 356698 640500 356704 640512
rect 356756 640500 356762 640552
rect 357894 640500 357900 640552
rect 357952 640540 357958 640552
rect 396534 640540 396540 640552
rect 357952 640512 396540 640540
rect 357952 640500 357958 640512
rect 396534 640500 396540 640512
rect 396592 640500 396598 640552
rect 315206 640432 315212 640484
rect 315264 640472 315270 640484
rect 322382 640472 322388 640484
rect 315264 640444 322388 640472
rect 315264 640432 315270 640444
rect 322382 640432 322388 640444
rect 322440 640432 322446 640484
rect 360010 640432 360016 640484
rect 360068 640472 360074 640484
rect 379422 640472 379428 640484
rect 360068 640444 379428 640472
rect 360068 640432 360074 640444
rect 379422 640432 379428 640444
rect 379480 640432 379486 640484
rect 310330 640364 310336 640416
rect 310388 640404 310394 640416
rect 320818 640404 320824 640416
rect 310388 640376 320824 640404
rect 310388 640364 310394 640376
rect 320818 640364 320824 640376
rect 320876 640364 320882 640416
rect 361206 640364 361212 640416
rect 361264 640404 361270 640416
rect 384390 640404 384396 640416
rect 361264 640376 384396 640404
rect 361264 640364 361270 640376
rect 384390 640364 384396 640376
rect 384448 640364 384454 640416
rect 254486 640296 254492 640348
rect 254544 640336 254550 640348
rect 273990 640336 273996 640348
rect 254544 640308 273996 640336
rect 254544 640296 254550 640308
rect 273990 640296 273996 640308
rect 274048 640296 274054 640348
rect 311802 640296 311808 640348
rect 311860 640336 311866 640348
rect 323578 640336 323584 640348
rect 311860 640308 323584 640336
rect 311860 640296 311866 640308
rect 323578 640296 323584 640308
rect 323636 640296 323642 640348
rect 361114 640296 361120 640348
rect 361172 640336 361178 640348
rect 385494 640336 385500 640348
rect 361172 640308 385500 640336
rect 361172 640296 361178 640308
rect 385494 640296 385500 640308
rect 385552 640296 385558 640348
rect 367554 639956 367560 640008
rect 367612 639996 367618 640008
rect 367612 639968 389174 639996
rect 367612 639956 367618 639968
rect 364794 639888 364800 639940
rect 364852 639928 364858 639940
rect 373258 639928 373264 639940
rect 364852 639900 373264 639928
rect 364852 639888 364858 639900
rect 373258 639888 373264 639900
rect 373316 639888 373322 639940
rect 365714 639820 365720 639872
rect 365772 639860 365778 639872
rect 373166 639860 373172 639872
rect 365772 639832 373172 639860
rect 365772 639820 365778 639832
rect 373166 639820 373172 639832
rect 373224 639820 373230 639872
rect 368106 639752 368112 639804
rect 368164 639792 368170 639804
rect 372338 639792 372344 639804
rect 368164 639764 372344 639792
rect 368164 639752 368170 639764
rect 372338 639752 372344 639764
rect 372396 639752 372402 639804
rect 327718 639684 327724 639736
rect 327776 639724 327782 639736
rect 382366 639724 382372 639736
rect 327776 639696 382372 639724
rect 327776 639684 327782 639696
rect 382366 639684 382372 639696
rect 382424 639684 382430 639736
rect 358446 639616 358452 639668
rect 358504 639656 358510 639668
rect 374638 639656 374644 639668
rect 358504 639628 374644 639656
rect 358504 639616 358510 639628
rect 374638 639616 374644 639628
rect 374696 639616 374702 639668
rect 377490 639616 377496 639668
rect 377548 639656 377554 639668
rect 377548 639628 385816 639656
rect 377548 639616 377554 639628
rect 358630 639548 358636 639600
rect 358688 639588 358694 639600
rect 376294 639588 376300 639600
rect 358688 639560 376300 639588
rect 358688 639548 358694 639560
rect 376294 639548 376300 639560
rect 376352 639548 376358 639600
rect 385678 639588 385684 639600
rect 381556 639560 385684 639588
rect 319714 639480 319720 639532
rect 319772 639520 319778 639532
rect 378502 639520 378508 639532
rect 319772 639492 378508 639520
rect 319772 639480 319778 639492
rect 378502 639480 378508 639492
rect 378560 639480 378566 639532
rect 319530 639412 319536 639464
rect 319588 639452 319594 639464
rect 380158 639452 380164 639464
rect 319588 639424 380164 639452
rect 319588 639412 319594 639424
rect 380158 639412 380164 639424
rect 380216 639412 380222 639464
rect 319162 639344 319168 639396
rect 319220 639384 319226 639396
rect 322474 639384 322480 639396
rect 319220 639356 322480 639384
rect 319220 639344 319226 639356
rect 322474 639344 322480 639356
rect 322532 639344 322538 639396
rect 358906 639344 358912 639396
rect 358964 639384 358970 639396
rect 371878 639384 371884 639396
rect 358964 639356 371884 639384
rect 358964 639344 358970 639356
rect 371878 639344 371884 639356
rect 371936 639344 371942 639396
rect 372338 639344 372344 639396
rect 372396 639344 372402 639396
rect 373074 639344 373080 639396
rect 373132 639344 373138 639396
rect 373166 639344 373172 639396
rect 373224 639344 373230 639396
rect 373258 639344 373264 639396
rect 373316 639344 373322 639396
rect 373994 639344 374000 639396
rect 374052 639344 374058 639396
rect 381262 639384 381268 639396
rect 376726 639356 381268 639384
rect 292022 639276 292028 639328
rect 292080 639276 292086 639328
rect 294046 639276 294052 639328
rect 294104 639316 294110 639328
rect 294104 639288 296714 639316
rect 294104 639276 294110 639288
rect 292040 638976 292068 639276
rect 296686 639112 296714 639288
rect 305086 639276 305092 639328
rect 305144 639316 305150 639328
rect 305144 639288 306374 639316
rect 305144 639276 305150 639288
rect 306346 639180 306374 639288
rect 307478 639276 307484 639328
rect 307536 639276 307542 639328
rect 309686 639276 309692 639328
rect 309744 639316 309750 639328
rect 354030 639316 354036 639328
rect 309744 639288 354036 639316
rect 309744 639276 309750 639288
rect 354030 639276 354036 639288
rect 354088 639276 354094 639328
rect 370590 639276 370596 639328
rect 370648 639276 370654 639328
rect 307496 639248 307524 639276
rect 351270 639248 351276 639260
rect 307496 639220 351276 639248
rect 351270 639208 351276 639220
rect 351328 639208 351334 639260
rect 353938 639180 353944 639192
rect 306346 639152 353944 639180
rect 353938 639140 353944 639152
rect 353996 639140 354002 639192
rect 322198 639112 322204 639124
rect 296686 639084 322204 639112
rect 322198 639072 322204 639084
rect 322256 639072 322262 639124
rect 361482 639004 361488 639056
rect 361540 639044 361546 639056
rect 370608 639044 370636 639276
rect 361540 639016 370636 639044
rect 361540 639004 361546 639016
rect 322290 638976 322296 638988
rect 292040 638948 322296 638976
rect 322290 638936 322296 638948
rect 322348 638936 322354 638988
rect 372356 638976 372384 639344
rect 373092 639044 373120 639344
rect 373184 639180 373212 639344
rect 373276 639248 373304 639344
rect 374012 639316 374040 639344
rect 376726 639316 376754 639356
rect 381262 639344 381268 639356
rect 381320 639344 381326 639396
rect 374012 639288 376754 639316
rect 381556 639248 381584 639560
rect 385678 639548 385684 639560
rect 385736 639548 385742 639600
rect 381722 639344 381728 639396
rect 381780 639344 381786 639396
rect 373276 639220 381584 639248
rect 381740 639180 381768 639344
rect 373184 639152 381768 639180
rect 385788 639112 385816 639628
rect 389146 639588 389174 639968
rect 401778 639588 401784 639600
rect 389146 639560 401784 639588
rect 401778 639548 401784 639560
rect 401836 639548 401842 639600
rect 396258 639412 396264 639464
rect 396316 639452 396322 639464
rect 399018 639452 399024 639464
rect 396316 639424 399024 639452
rect 396316 639412 396322 639424
rect 399018 639412 399024 639424
rect 399076 639412 399082 639464
rect 385862 639344 385868 639396
rect 385920 639344 385926 639396
rect 385954 639344 385960 639396
rect 386012 639384 386018 639396
rect 386012 639356 386092 639384
rect 386012 639344 386018 639356
rect 385880 639180 385908 639344
rect 386064 639248 386092 639356
rect 386138 639344 386144 639396
rect 386196 639344 386202 639396
rect 397914 639344 397920 639396
rect 397972 639384 397978 639396
rect 398834 639384 398840 639396
rect 397972 639356 398840 639384
rect 397972 639344 397978 639356
rect 398834 639344 398840 639356
rect 398892 639344 398898 639396
rect 386156 639316 386184 639344
rect 400214 639316 400220 639328
rect 386156 639288 400220 639316
rect 400214 639276 400220 639288
rect 400272 639276 400278 639328
rect 402330 639248 402336 639260
rect 386064 639220 402336 639248
rect 402330 639208 402336 639220
rect 402388 639208 402394 639260
rect 401962 639180 401968 639192
rect 385880 639152 401968 639180
rect 401962 639140 401968 639152
rect 402020 639140 402026 639192
rect 400398 639112 400404 639124
rect 385788 639084 400404 639112
rect 400398 639072 400404 639084
rect 400456 639072 400462 639124
rect 402514 639044 402520 639056
rect 373092 639016 381492 639044
rect 372356 638948 376754 638976
rect 376726 638840 376754 638948
rect 381464 638908 381492 639016
rect 384868 639016 402520 639044
rect 384868 638908 384896 639016
rect 402514 639004 402520 639016
rect 402572 639004 402578 639056
rect 403894 638976 403900 638988
rect 381464 638880 384896 638908
rect 384960 638948 403900 638976
rect 384960 638840 384988 638948
rect 403894 638936 403900 638948
rect 403952 638936 403958 638988
rect 376726 638812 384988 638840
rect 49418 636692 49424 636744
rect 49476 636732 49482 636744
rect 50522 636732 50528 636744
rect 49476 636704 50528 636732
rect 49476 636692 49482 636704
rect 50522 636692 50528 636704
rect 50580 636692 50586 636744
rect 403618 634788 403624 634840
rect 403676 634828 403682 634840
rect 478690 634828 478696 634840
rect 403676 634800 478696 634828
rect 403676 634788 403682 634800
rect 478690 634788 478696 634800
rect 478748 634788 478754 634840
rect 254394 633428 254400 633480
rect 254452 633468 254458 633480
rect 271230 633468 271236 633480
rect 254452 633440 271236 633468
rect 254452 633428 254458 633440
rect 271230 633428 271236 633440
rect 271288 633428 271294 633480
rect 523678 632000 523684 632052
rect 523736 632040 523742 632052
rect 580166 632040 580172 632052
rect 523736 632012 580172 632040
rect 523736 632000 523742 632012
rect 580166 632000 580172 632012
rect 580224 632000 580230 632052
rect 49142 629348 49148 629400
rect 49200 629388 49206 629400
rect 50430 629388 50436 629400
rect 49200 629360 50436 629388
rect 49200 629348 49206 629360
rect 50430 629348 50436 629360
rect 50488 629348 50494 629400
rect 254302 627920 254308 627972
rect 254360 627960 254366 627972
rect 278038 627960 278044 627972
rect 254360 627932 278044 627960
rect 254360 627920 254366 627932
rect 278038 627920 278044 627932
rect 278096 627920 278102 627972
rect 254026 622412 254032 622464
rect 254084 622452 254090 622464
rect 264238 622452 264244 622464
rect 254084 622424 264244 622452
rect 254084 622412 254090 622424
rect 264238 622412 264244 622424
rect 264296 622412 264302 622464
rect 48774 619012 48780 619064
rect 48832 619052 48838 619064
rect 50338 619052 50344 619064
rect 48832 619024 50344 619052
rect 48832 619012 48838 619024
rect 50338 619012 50344 619024
rect 50396 619012 50402 619064
rect 538858 616836 538864 616888
rect 538916 616876 538922 616888
rect 580166 616876 580172 616888
rect 538916 616848 580172 616876
rect 538916 616836 538922 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 254486 611328 254492 611380
rect 254544 611368 254550 611380
rect 269758 611368 269764 611380
rect 254544 611340 269764 611368
rect 254544 611328 254550 611340
rect 269758 611328 269764 611340
rect 269816 611328 269822 611380
rect 254210 604460 254216 604512
rect 254268 604500 254274 604512
rect 275278 604500 275284 604512
rect 254268 604472 275284 604500
rect 254268 604460 254274 604472
rect 275278 604460 275284 604472
rect 275336 604460 275342 604512
rect 398374 600244 398380 600296
rect 398432 600284 398438 600296
rect 403618 600284 403624 600296
rect 398432 600256 403624 600284
rect 398432 600244 398438 600256
rect 403618 600244 403624 600256
rect 403676 600244 403682 600296
rect 364794 600176 364800 600228
rect 364852 600216 364858 600228
rect 365162 600216 365168 600228
rect 364852 600188 365168 600216
rect 364852 600176 364858 600188
rect 365162 600176 365168 600188
rect 365220 600176 365226 600228
rect 300946 599836 300952 599888
rect 301004 599876 301010 599888
rect 302188 599876 302194 599888
rect 301004 599848 302194 599876
rect 301004 599836 301010 599848
rect 302188 599836 302194 599848
rect 302246 599836 302252 599888
rect 306374 599836 306380 599888
rect 306432 599876 306438 599888
rect 307708 599876 307714 599888
rect 306432 599848 307714 599876
rect 306432 599836 306438 599848
rect 307708 599836 307714 599848
rect 307766 599836 307772 599888
rect 382274 599836 382280 599888
rect 382332 599876 382338 599888
rect 400582 599876 400588 599888
rect 382332 599848 400588 599876
rect 382332 599836 382338 599848
rect 400582 599836 400588 599848
rect 400640 599836 400646 599888
rect 379790 599768 379796 599820
rect 379848 599808 379854 599820
rect 399202 599808 399208 599820
rect 379848 599780 399208 599808
rect 379848 599768 379854 599780
rect 399202 599768 399208 599780
rect 399260 599768 399266 599820
rect 378410 599700 378416 599752
rect 378468 599740 378474 599752
rect 399294 599740 399300 599752
rect 378468 599712 399300 599740
rect 378468 599700 378474 599712
rect 399294 599700 399300 599712
rect 399352 599700 399358 599752
rect 372614 599632 372620 599684
rect 372672 599672 372678 599684
rect 399386 599672 399392 599684
rect 372672 599644 399392 599672
rect 372672 599632 372678 599644
rect 399386 599632 399392 599644
rect 399444 599632 399450 599684
rect 365714 599564 365720 599616
rect 365772 599604 365778 599616
rect 400490 599604 400496 599616
rect 365772 599576 400496 599604
rect 365772 599564 365778 599576
rect 400490 599564 400496 599576
rect 400548 599564 400554 599616
rect 300854 599360 300860 599412
rect 300912 599400 300918 599412
rect 301406 599400 301412 599412
rect 300912 599372 301412 599400
rect 300912 599360 300918 599372
rect 301406 599360 301412 599372
rect 301464 599400 301470 599412
rect 357066 599400 357072 599412
rect 301464 599372 357072 599400
rect 301464 599360 301470 599372
rect 357066 599360 357072 599372
rect 357124 599360 357130 599412
rect 283006 599292 283012 599344
rect 283064 599332 283070 599344
rect 333238 599332 333244 599344
rect 283064 599304 333244 599332
rect 283064 599292 283070 599304
rect 333238 599292 333244 599304
rect 333296 599292 333302 599344
rect 304994 599224 305000 599276
rect 305052 599264 305058 599276
rect 305914 599264 305920 599276
rect 305052 599236 305920 599264
rect 305052 599224 305058 599236
rect 305914 599224 305920 599236
rect 305972 599264 305978 599276
rect 355594 599264 355600 599276
rect 305972 599236 355600 599264
rect 305972 599224 305978 599236
rect 355594 599224 355600 599236
rect 355652 599224 355658 599276
rect 302142 599156 302148 599208
rect 302200 599196 302206 599208
rect 353202 599196 353208 599208
rect 302200 599168 353208 599196
rect 302200 599156 302206 599168
rect 353202 599156 353208 599168
rect 353260 599156 353266 599208
rect 359642 599156 359648 599208
rect 359700 599196 359706 599208
rect 360010 599196 360016 599208
rect 359700 599168 360016 599196
rect 359700 599156 359706 599168
rect 360010 599156 360016 599168
rect 360068 599196 360074 599208
rect 404722 599196 404728 599208
rect 360068 599168 404728 599196
rect 360068 599156 360074 599168
rect 404722 599156 404728 599168
rect 404780 599156 404786 599208
rect 296714 599088 296720 599140
rect 296772 599128 296778 599140
rect 298002 599128 298008 599140
rect 296772 599100 298008 599128
rect 296772 599088 296778 599100
rect 298002 599088 298008 599100
rect 298060 599128 298066 599140
rect 349890 599128 349896 599140
rect 298060 599100 349896 599128
rect 298060 599088 298066 599100
rect 349890 599088 349896 599100
rect 349948 599088 349954 599140
rect 387702 599088 387708 599140
rect 387760 599128 387766 599140
rect 404998 599128 405004 599140
rect 387760 599100 405004 599128
rect 387760 599088 387766 599100
rect 404998 599088 405004 599100
rect 405056 599088 405062 599140
rect 353110 599020 353116 599072
rect 353168 599060 353174 599072
rect 361574 599060 361580 599072
rect 353168 599032 361580 599060
rect 353168 599020 353174 599032
rect 361574 599020 361580 599032
rect 361632 599060 361638 599072
rect 361758 599060 361764 599072
rect 361632 599032 361764 599060
rect 361632 599020 361638 599032
rect 361758 599020 361764 599032
rect 361816 599060 361822 599072
rect 472618 599060 472624 599072
rect 361816 599032 472624 599060
rect 361816 599020 361822 599032
rect 472618 599020 472624 599032
rect 472676 599020 472682 599072
rect 254118 598952 254124 599004
rect 254176 598992 254182 599004
rect 273898 598992 273904 599004
rect 254176 598964 273904 598992
rect 254176 598952 254182 598964
rect 273898 598952 273904 598964
rect 273956 598952 273962 599004
rect 299474 598952 299480 599004
rect 299532 598992 299538 599004
rect 300302 598992 300308 599004
rect 299532 598964 300308 598992
rect 299532 598952 299538 598964
rect 300302 598952 300308 598964
rect 300360 598992 300366 599004
rect 361022 598992 361028 599004
rect 300360 598964 361028 598992
rect 300360 598952 300366 598964
rect 361022 598952 361028 598964
rect 361080 598952 361086 599004
rect 386598 598952 386604 599004
rect 386656 598992 386662 599004
rect 387702 598992 387708 599004
rect 386656 598964 387708 598992
rect 386656 598952 386662 598964
rect 387702 598952 387708 598964
rect 387760 598952 387766 599004
rect 299382 598884 299388 598936
rect 299440 598924 299446 598936
rect 359642 598924 359648 598936
rect 299440 598896 359648 598924
rect 299440 598884 299446 598896
rect 359642 598884 359648 598896
rect 359700 598884 359706 598936
rect 388254 598884 388260 598936
rect 388312 598924 388318 598936
rect 521746 598924 521752 598936
rect 388312 598896 521752 598924
rect 388312 598884 388318 598896
rect 521746 598884 521752 598896
rect 521804 598884 521810 598936
rect 304718 598816 304724 598868
rect 304776 598856 304782 598868
rect 361206 598856 361212 598868
rect 304776 598828 361212 598856
rect 304776 598816 304782 598828
rect 361206 598816 361212 598828
rect 361264 598816 361270 598868
rect 386414 598816 386420 598868
rect 386472 598856 386478 598868
rect 387150 598856 387156 598868
rect 386472 598828 387156 598856
rect 386472 598816 386478 598828
rect 387150 598816 387156 598828
rect 387208 598856 387214 598868
rect 513834 598856 513840 598868
rect 387208 598828 513840 598856
rect 387208 598816 387214 598828
rect 513834 598816 513840 598828
rect 513892 598816 513898 598868
rect 298646 598748 298652 598800
rect 298704 598788 298710 598800
rect 299382 598788 299388 598800
rect 298704 598760 299388 598788
rect 298704 598748 298710 598760
rect 299382 598748 299388 598760
rect 299440 598788 299446 598800
rect 355502 598788 355508 598800
rect 299440 598760 355508 598788
rect 299440 598748 299446 598760
rect 355502 598748 355508 598760
rect 355560 598748 355566 598800
rect 388438 598748 388444 598800
rect 388496 598788 388502 598800
rect 478138 598788 478144 598800
rect 388496 598760 478144 598788
rect 388496 598748 388502 598760
rect 478138 598748 478144 598760
rect 478196 598748 478202 598800
rect 305822 598680 305828 598732
rect 305880 598720 305886 598732
rect 306282 598720 306288 598732
rect 305880 598692 306288 598720
rect 305880 598680 305886 598692
rect 306282 598680 306288 598692
rect 306340 598720 306346 598732
rect 361114 598720 361120 598732
rect 306340 598692 361120 598720
rect 306340 598680 306346 598692
rect 361114 598680 361120 598692
rect 361172 598680 361178 598732
rect 304166 598612 304172 598664
rect 304224 598652 304230 598664
rect 304626 598652 304632 598664
rect 304224 598624 304632 598652
rect 304224 598612 304230 598624
rect 304626 598612 304632 598624
rect 304684 598652 304690 598664
rect 357158 598652 357164 598664
rect 304684 598624 357164 598652
rect 304684 598612 304690 598624
rect 357158 598612 357164 598624
rect 357216 598612 357222 598664
rect 361022 598612 361028 598664
rect 361080 598652 361086 598664
rect 381078 598652 381084 598664
rect 361080 598624 381084 598652
rect 361080 598612 361086 598624
rect 381078 598612 381084 598624
rect 381136 598612 381142 598664
rect 304902 598544 304908 598596
rect 304960 598584 304966 598596
rect 342898 598584 342904 598596
rect 304960 598556 342904 598584
rect 304960 598544 304966 598556
rect 342898 598544 342904 598556
rect 342956 598544 342962 598596
rect 363598 598544 363604 598596
rect 363656 598584 363662 598596
rect 371694 598584 371700 598596
rect 363656 598556 371700 598584
rect 363656 598544 363662 598556
rect 371694 598544 371700 598556
rect 371752 598544 371758 598596
rect 377214 598544 377220 598596
rect 377272 598584 377278 598596
rect 397638 598584 397644 598596
rect 377272 598556 397644 598584
rect 377272 598544 377278 598556
rect 397638 598544 397644 598556
rect 397696 598544 397702 598596
rect 294506 598476 294512 598528
rect 294564 598516 294570 598528
rect 300118 598516 300124 598528
rect 294564 598488 300124 598516
rect 294564 598476 294570 598488
rect 300118 598476 300124 598488
rect 300176 598476 300182 598528
rect 308306 598476 308312 598528
rect 308364 598516 308370 598528
rect 357066 598516 357072 598528
rect 308364 598488 357072 598516
rect 308364 598476 308370 598488
rect 357066 598476 357072 598488
rect 357124 598476 357130 598528
rect 366174 598476 366180 598528
rect 366232 598516 366238 598528
rect 397730 598516 397736 598528
rect 366232 598488 397736 598516
rect 366232 598476 366238 598488
rect 397730 598476 397736 598488
rect 397788 598476 397794 598528
rect 317322 598408 317328 598460
rect 317380 598448 317386 598460
rect 401042 598448 401048 598460
rect 317380 598420 401048 598448
rect 317380 598408 317386 598420
rect 401042 598408 401048 598420
rect 401100 598408 401106 598460
rect 290918 598340 290924 598392
rect 290976 598380 290982 598392
rect 404630 598380 404636 598392
rect 290976 598352 404636 598380
rect 290976 598340 290982 598352
rect 404630 598340 404636 598352
rect 404688 598340 404694 598392
rect 288986 598272 288992 598324
rect 289044 598312 289050 598324
rect 403250 598312 403256 598324
rect 289044 598284 403256 598312
rect 289044 598272 289050 598284
rect 403250 598272 403256 598284
rect 403308 598272 403314 598324
rect 284570 598204 284576 598256
rect 284628 598244 284634 598256
rect 403342 598244 403348 598256
rect 284628 598216 403348 598244
rect 284628 598204 284634 598216
rect 403342 598204 403348 598216
rect 403400 598204 403406 598256
rect 471238 598204 471244 598256
rect 471296 598244 471302 598256
rect 496446 598244 496452 598256
rect 471296 598216 496452 598244
rect 471296 598204 471302 598216
rect 496446 598204 496452 598216
rect 496504 598204 496510 598256
rect 282914 598136 282920 598188
rect 282972 598176 282978 598188
rect 283650 598176 283656 598188
rect 282972 598148 283656 598176
rect 282972 598136 282978 598148
rect 283650 598136 283656 598148
rect 283708 598136 283714 598188
rect 285582 598136 285588 598188
rect 285640 598176 285646 598188
rect 286318 598176 286324 598188
rect 285640 598148 286324 598176
rect 285640 598136 285646 598148
rect 286318 598136 286324 598148
rect 286376 598136 286382 598188
rect 291102 598136 291108 598188
rect 291160 598176 291166 598188
rect 291838 598176 291844 598188
rect 291160 598148 291844 598176
rect 291160 598136 291166 598148
rect 291838 598136 291844 598148
rect 291896 598136 291902 598188
rect 292574 598136 292580 598188
rect 292632 598176 292638 598188
rect 293586 598176 293592 598188
rect 292632 598148 293592 598176
rect 292632 598136 292638 598148
rect 293586 598136 293592 598148
rect 293644 598136 293650 598188
rect 295334 598136 295340 598188
rect 295392 598176 295398 598188
rect 295794 598176 295800 598188
rect 295392 598148 295800 598176
rect 295392 598136 295398 598148
rect 295794 598136 295800 598148
rect 295852 598136 295858 598188
rect 299198 598136 299204 598188
rect 299256 598176 299262 598188
rect 300670 598176 300676 598188
rect 299256 598148 300676 598176
rect 299256 598136 299262 598148
rect 300670 598136 300676 598148
rect 300728 598136 300734 598188
rect 302878 598136 302884 598188
rect 302936 598176 302942 598188
rect 311066 598176 311072 598188
rect 302936 598148 311072 598176
rect 302936 598136 302942 598148
rect 311066 598136 311072 598148
rect 311124 598136 311130 598188
rect 311986 598136 311992 598188
rect 312044 598176 312050 598188
rect 312906 598176 312912 598188
rect 312044 598148 312912 598176
rect 312044 598136 312050 598148
rect 312906 598136 312912 598148
rect 312964 598136 312970 598188
rect 313274 598136 313280 598188
rect 313332 598176 313338 598188
rect 314010 598176 314016 598188
rect 313332 598148 314016 598176
rect 313332 598136 313338 598148
rect 314010 598136 314016 598148
rect 314068 598136 314074 598188
rect 314654 598136 314660 598188
rect 314712 598176 314718 598188
rect 315114 598176 315120 598188
rect 314712 598148 315120 598176
rect 314712 598136 314718 598148
rect 315114 598136 315120 598148
rect 315172 598136 315178 598188
rect 316862 598136 316868 598188
rect 316920 598176 316926 598188
rect 324958 598176 324964 598188
rect 316920 598148 324964 598176
rect 316920 598136 316926 598148
rect 324958 598136 324964 598148
rect 325016 598136 325022 598188
rect 364426 598136 364432 598188
rect 364484 598176 364490 598188
rect 365254 598176 365260 598188
rect 364484 598148 365260 598176
rect 364484 598136 364490 598148
rect 365254 598136 365260 598148
rect 365312 598136 365318 598188
rect 367094 598136 367100 598188
rect 367152 598176 367158 598188
rect 368014 598176 368020 598188
rect 367152 598148 368020 598176
rect 367152 598136 367158 598148
rect 368014 598136 368020 598148
rect 368072 598136 368078 598188
rect 372798 598136 372804 598188
rect 372856 598176 372862 598188
rect 372982 598176 372988 598188
rect 372856 598148 372988 598176
rect 372856 598136 372862 598148
rect 372982 598136 372988 598148
rect 373040 598136 373046 598188
rect 376662 598136 376668 598188
rect 376720 598176 376726 598188
rect 377398 598176 377404 598188
rect 376720 598148 377404 598176
rect 376720 598136 376726 598148
rect 377398 598136 377404 598148
rect 377456 598136 377462 598188
rect 378318 598136 378324 598188
rect 378376 598176 378382 598188
rect 379054 598176 379060 598188
rect 378376 598148 379060 598176
rect 378376 598136 378382 598148
rect 379054 598136 379060 598148
rect 379112 598136 379118 598188
rect 379606 598136 379612 598188
rect 379664 598176 379670 598188
rect 380158 598176 380164 598188
rect 379664 598148 380164 598176
rect 379664 598136 379670 598148
rect 380158 598136 380164 598148
rect 380216 598136 380222 598188
rect 380986 598136 380992 598188
rect 381044 598176 381050 598188
rect 381814 598176 381820 598188
rect 381044 598148 381820 598176
rect 381044 598136 381050 598148
rect 381814 598136 381820 598148
rect 381872 598136 381878 598188
rect 382366 598136 382372 598188
rect 382424 598176 382430 598188
rect 382918 598176 382924 598188
rect 382424 598148 382924 598176
rect 382424 598136 382430 598148
rect 382918 598136 382924 598148
rect 382976 598136 382982 598188
rect 385034 598136 385040 598188
rect 385092 598176 385098 598188
rect 385678 598176 385684 598188
rect 385092 598148 385684 598176
rect 385092 598136 385098 598148
rect 385678 598136 385684 598148
rect 385736 598136 385742 598188
rect 388254 598136 388260 598188
rect 388312 598176 388318 598188
rect 388530 598176 388536 598188
rect 388312 598148 388536 598176
rect 388312 598136 388318 598148
rect 388530 598136 388536 598148
rect 388588 598136 388594 598188
rect 389266 598136 389272 598188
rect 389324 598176 389330 598188
rect 390094 598176 390100 598188
rect 389324 598148 390100 598176
rect 389324 598136 389330 598148
rect 390094 598136 390100 598148
rect 390152 598136 390158 598188
rect 393314 598136 393320 598188
rect 393372 598176 393378 598188
rect 393958 598176 393964 598188
rect 393372 598148 393964 598176
rect 393372 598136 393378 598148
rect 393958 598136 393964 598148
rect 394016 598136 394022 598188
rect 394694 598136 394700 598188
rect 394752 598176 394758 598188
rect 395062 598176 395068 598188
rect 394752 598148 395068 598176
rect 394752 598136 394758 598148
rect 395062 598136 395068 598148
rect 395120 598136 395126 598188
rect 396074 598136 396080 598188
rect 396132 598176 396138 598188
rect 396718 598176 396724 598188
rect 396132 598148 396724 598176
rect 396132 598136 396138 598148
rect 396718 598136 396724 598148
rect 396776 598136 396782 598188
rect 291194 598068 291200 598120
rect 291252 598108 291258 598120
rect 291930 598108 291936 598120
rect 291252 598080 291936 598108
rect 291252 598068 291258 598080
rect 291930 598068 291936 598080
rect 291988 598068 291994 598120
rect 309134 598068 309140 598120
rect 309192 598108 309198 598120
rect 310146 598108 310152 598120
rect 309192 598080 310152 598108
rect 309192 598068 309198 598080
rect 310146 598068 310152 598080
rect 310204 598068 310210 598120
rect 311894 598068 311900 598120
rect 311952 598108 311958 598120
rect 312354 598108 312360 598120
rect 311952 598080 312360 598108
rect 311952 598068 311958 598080
rect 312354 598068 312360 598080
rect 312412 598068 312418 598120
rect 372706 598068 372712 598120
rect 372764 598108 372770 598120
rect 373534 598108 373540 598120
rect 372764 598080 373540 598108
rect 372764 598068 372770 598080
rect 373534 598068 373540 598080
rect 373592 598068 373598 598120
rect 300762 598000 300768 598052
rect 300820 598040 300826 598052
rect 319530 598040 319536 598052
rect 300820 598012 319536 598040
rect 300820 598000 300826 598012
rect 319530 598000 319536 598012
rect 319588 598000 319594 598052
rect 290366 597796 290372 597848
rect 290424 597836 290430 597848
rect 294598 597836 294604 597848
rect 290424 597808 294604 597836
rect 290424 597796 290430 597808
rect 294598 597796 294604 597808
rect 294656 597796 294662 597848
rect 286870 597592 286876 597644
rect 286928 597632 286934 597644
rect 289078 597632 289084 597644
rect 286928 597604 289084 597632
rect 286928 597592 286934 597604
rect 289078 597592 289084 597604
rect 289136 597592 289142 597644
rect 390554 597592 390560 597644
rect 390612 597632 390618 597644
rect 391198 597632 391204 597644
rect 390612 597604 391204 597632
rect 390612 597592 390618 597604
rect 391198 597592 391204 597604
rect 391256 597592 391262 597644
rect 327718 596912 327724 596964
rect 327776 596912 327782 596964
rect 311066 596844 311072 596896
rect 311124 596884 311130 596896
rect 327736 596884 327764 596912
rect 335998 596884 336004 596896
rect 311124 596856 336004 596884
rect 311124 596844 311130 596856
rect 335998 596844 336004 596856
rect 336056 596844 336062 596896
rect 342162 596844 342168 596896
rect 342220 596884 342226 596896
rect 363966 596884 363972 596896
rect 342220 596856 363972 596884
rect 342220 596844 342226 596856
rect 363966 596844 363972 596856
rect 364024 596844 364030 596896
rect 297542 596776 297548 596828
rect 297600 596816 297606 596828
rect 327718 596816 327724 596828
rect 297600 596788 327724 596816
rect 297600 596776 297606 596788
rect 327718 596776 327724 596788
rect 327776 596776 327782 596828
rect 329098 596776 329104 596828
rect 329156 596816 329162 596828
rect 398190 596816 398196 596828
rect 329156 596788 398196 596816
rect 329156 596776 329162 596788
rect 398190 596776 398196 596788
rect 398248 596776 398254 596828
rect 384390 596572 384396 596624
rect 384448 596612 384454 596624
rect 392578 596612 392584 596624
rect 384448 596584 392584 596612
rect 384448 596572 384454 596584
rect 392578 596572 392584 596584
rect 392636 596572 392642 596624
rect 302234 595552 302240 595604
rect 302292 595592 302298 595604
rect 334618 595592 334624 595604
rect 302292 595564 334624 595592
rect 302292 595552 302298 595564
rect 334618 595552 334624 595564
rect 334676 595552 334682 595604
rect 362954 595552 362960 595604
rect 363012 595592 363018 595604
rect 387794 595592 387800 595604
rect 363012 595564 387800 595592
rect 363012 595552 363018 595564
rect 387794 595552 387800 595564
rect 387852 595552 387858 595604
rect 333882 595484 333888 595536
rect 333940 595524 333946 595536
rect 367370 595524 367376 595536
rect 333940 595496 367376 595524
rect 333940 595484 333946 595496
rect 367370 595484 367376 595496
rect 367428 595484 367434 595536
rect 291286 595416 291292 595468
rect 291344 595456 291350 595468
rect 345658 595456 345664 595468
rect 291344 595428 345664 595456
rect 291344 595416 291350 595428
rect 345658 595416 345664 595428
rect 345716 595416 345722 595468
rect 347774 595416 347780 595468
rect 347832 595456 347838 595468
rect 510706 595456 510712 595468
rect 347832 595428 510712 595456
rect 347832 595416 347838 595428
rect 510706 595416 510712 595428
rect 510764 595416 510770 595468
rect 49510 594804 49516 594856
rect 49568 594844 49574 594856
rect 51810 594844 51816 594856
rect 49568 594816 51816 594844
rect 49568 594804 49574 594816
rect 51810 594804 51816 594816
rect 51868 594804 51874 594856
rect 288066 594192 288072 594244
rect 288124 594232 288130 594244
rect 331950 594232 331956 594244
rect 288124 594204 331956 594232
rect 288124 594192 288130 594204
rect 331950 594192 331956 594204
rect 332008 594192 332014 594244
rect 324222 594124 324228 594176
rect 324280 594164 324286 594176
rect 375374 594164 375380 594176
rect 324280 594136 375380 594164
rect 324280 594124 324286 594136
rect 375374 594124 375380 594136
rect 375432 594124 375438 594176
rect 381538 594124 381544 594176
rect 381596 594164 381602 594176
rect 386414 594164 386420 594176
rect 381596 594136 386420 594164
rect 381596 594124 381602 594136
rect 386414 594124 386420 594136
rect 386472 594124 386478 594176
rect 311158 594056 311164 594108
rect 311216 594096 311222 594108
rect 327810 594096 327816 594108
rect 311216 594068 327816 594096
rect 311216 594056 311222 594068
rect 327810 594056 327816 594068
rect 327868 594056 327874 594108
rect 331214 594056 331220 594108
rect 331272 594096 331278 594108
rect 499574 594096 499580 594108
rect 331272 594068 499580 594096
rect 331272 594056 331278 594068
rect 499574 594056 499580 594068
rect 499632 594056 499638 594108
rect 254762 593376 254768 593428
rect 254820 593416 254826 593428
rect 271138 593416 271144 593428
rect 254820 593388 271144 593416
rect 254820 593376 254826 593388
rect 271138 593376 271144 593388
rect 271196 593376 271202 593428
rect 266354 592628 266360 592680
rect 266412 592668 266418 592680
rect 498194 592668 498200 592680
rect 266412 592640 498200 592668
rect 266412 592628 266418 592640
rect 498194 592628 498200 592640
rect 498252 592628 498258 592680
rect 312078 591948 312084 592000
rect 312136 591988 312142 592000
rect 316678 591988 316684 592000
rect 312136 591960 316684 591988
rect 312136 591948 312142 591960
rect 316678 591948 316684 591960
rect 316736 591948 316742 592000
rect 325510 591336 325516 591388
rect 325568 591376 325574 591388
rect 364702 591376 364708 591388
rect 325568 591348 364708 591376
rect 325568 591336 325574 591348
rect 364702 591336 364708 591348
rect 364760 591336 364766 591388
rect 371878 591336 371884 591388
rect 371936 591376 371942 591388
rect 392026 591376 392032 591388
rect 371936 591348 392032 591376
rect 371936 591336 371942 591348
rect 392026 591336 392032 591348
rect 392084 591336 392090 591388
rect 293954 591268 293960 591320
rect 294012 591308 294018 591320
rect 386782 591308 386788 591320
rect 294012 591280 386788 591308
rect 294012 591268 294018 591280
rect 386782 591268 386788 591280
rect 386840 591268 386846 591320
rect 485866 590656 485872 590708
rect 485924 590696 485930 590708
rect 579798 590696 579804 590708
rect 485924 590668 579804 590696
rect 485924 590656 485930 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 49602 590588 49608 590640
rect 49660 590628 49666 590640
rect 51718 590628 51724 590640
rect 49660 590600 51724 590628
rect 49660 590588 49666 590600
rect 51718 590588 51724 590600
rect 51776 590588 51782 590640
rect 306742 589976 306748 590028
rect 306800 590016 306806 590028
rect 333238 590016 333244 590028
rect 306800 589988 333244 590016
rect 306800 589976 306806 589988
rect 333238 589976 333244 589988
rect 333296 589976 333302 590028
rect 336642 589976 336648 590028
rect 336700 590016 336706 590028
rect 369026 590016 369032 590028
rect 336700 589988 369032 590016
rect 336700 589976 336706 589988
rect 369026 589976 369032 589988
rect 369084 589976 369090 590028
rect 292942 589908 292948 589960
rect 293000 589948 293006 589960
rect 349890 589948 349896 589960
rect 293000 589920 349896 589948
rect 293000 589908 293006 589920
rect 349890 589908 349896 589920
rect 349948 589908 349954 589960
rect 361114 589908 361120 589960
rect 361172 589948 361178 589960
rect 391934 589948 391940 589960
rect 361172 589920 391940 589948
rect 361172 589908 361178 589920
rect 391934 589908 391940 589920
rect 391992 589908 391998 589960
rect 385678 589228 385684 589280
rect 385736 589268 385742 589280
rect 390646 589268 390652 589280
rect 385736 589240 390652 589268
rect 385736 589228 385742 589240
rect 390646 589228 390652 589240
rect 390704 589228 390710 589280
rect 311986 588616 311992 588668
rect 312044 588656 312050 588668
rect 338850 588656 338856 588668
rect 312044 588628 338856 588656
rect 312044 588616 312050 588628
rect 338850 588616 338856 588628
rect 338908 588616 338914 588668
rect 343542 588616 343548 588668
rect 343600 588656 343606 588668
rect 371786 588656 371792 588668
rect 343600 588628 371792 588656
rect 343600 588616 343606 588628
rect 371786 588616 371792 588628
rect 371844 588616 371850 588668
rect 288434 588548 288440 588600
rect 288492 588588 288498 588600
rect 347038 588588 347044 588600
rect 288492 588560 347044 588588
rect 288492 588548 288498 588560
rect 347038 588548 347044 588560
rect 347096 588548 347102 588600
rect 254486 587936 254492 587988
rect 254544 587976 254550 587988
rect 260098 587976 260104 587988
rect 254544 587948 260104 587976
rect 254544 587936 254550 587948
rect 260098 587936 260104 587948
rect 260156 587936 260162 587988
rect 329282 587120 329288 587172
rect 329340 587160 329346 587172
rect 372890 587160 372896 587172
rect 329340 587132 372896 587160
rect 329340 587120 329346 587132
rect 372890 587120 372896 587132
rect 372948 587120 372954 587172
rect 322474 585760 322480 585812
rect 322532 585800 322538 585812
rect 506474 585800 506480 585812
rect 322532 585772 506480 585800
rect 322532 585760 322538 585772
rect 506474 585760 506480 585772
rect 506532 585760 506538 585812
rect 340138 584536 340144 584588
rect 340196 584576 340202 584588
rect 396166 584576 396172 584588
rect 340196 584548 396172 584576
rect 340196 584536 340202 584548
rect 396166 584536 396172 584548
rect 396224 584536 396230 584588
rect 307754 584468 307760 584520
rect 307812 584508 307818 584520
rect 368566 584508 368572 584520
rect 307812 584480 368572 584508
rect 307812 584468 307818 584480
rect 368566 584468 368572 584480
rect 368624 584468 368630 584520
rect 287146 584400 287152 584452
rect 287204 584440 287210 584452
rect 353110 584440 353116 584452
rect 287204 584412 353116 584440
rect 287204 584400 287210 584412
rect 353110 584400 353116 584412
rect 353168 584400 353174 584452
rect 285674 582972 285680 583024
rect 285732 583012 285738 583024
rect 347130 583012 347136 583024
rect 285732 582984 347136 583012
rect 285732 582972 285738 582984
rect 347130 582972 347136 582984
rect 347188 582972 347194 583024
rect 385770 582360 385776 582412
rect 385828 582400 385834 582412
rect 389266 582400 389272 582412
rect 385828 582372 389272 582400
rect 385828 582360 385834 582372
rect 389266 582360 389272 582372
rect 389324 582360 389330 582412
rect 253934 581272 253940 581324
rect 253992 581312 253998 581324
rect 255958 581312 255964 581324
rect 253992 581284 255964 581312
rect 253992 581272 253998 581284
rect 255958 581272 255964 581284
rect 256016 581272 256022 581324
rect 310514 580252 310520 580304
rect 310572 580292 310578 580304
rect 374270 580292 374276 580304
rect 310572 580264 374276 580292
rect 310572 580252 310578 580264
rect 374270 580252 374276 580264
rect 374328 580252 374334 580304
rect 322382 578144 322388 578196
rect 322440 578184 322446 578196
rect 580166 578184 580172 578196
rect 322440 578156 580172 578184
rect 322440 578144 322446 578156
rect 580166 578144 580172 578156
rect 580224 578144 580230 578196
rect 300854 577464 300860 577516
rect 300912 577504 300918 577516
rect 342898 577504 342904 577516
rect 300912 577476 342904 577504
rect 300912 577464 300918 577476
rect 342898 577464 342904 577476
rect 342956 577464 342962 577516
rect 314838 576172 314844 576224
rect 314896 576212 314902 576224
rect 390646 576212 390652 576224
rect 314896 576184 390652 576212
rect 314896 576172 314902 576184
rect 390646 576172 390652 576184
rect 390704 576172 390710 576224
rect 286318 576104 286324 576156
rect 286376 576144 286382 576156
rect 386598 576144 386604 576156
rect 286376 576116 386604 576144
rect 286376 576104 286382 576116
rect 386598 576104 386604 576116
rect 386656 576104 386662 576156
rect 254486 575492 254492 575544
rect 254544 575532 254550 575544
rect 261478 575532 261484 575544
rect 254544 575504 261484 575532
rect 254544 575492 254550 575504
rect 261478 575492 261484 575504
rect 261536 575492 261542 575544
rect 323670 574744 323676 574796
rect 323728 574784 323734 574796
rect 382458 574784 382464 574796
rect 323728 574756 382464 574784
rect 323728 574744 323734 574756
rect 382458 574744 382464 574756
rect 382516 574744 382522 574796
rect 313366 573384 313372 573436
rect 313424 573424 313430 573436
rect 376938 573424 376944 573436
rect 313424 573396 376944 573424
rect 313424 573384 313430 573396
rect 376938 573384 376944 573396
rect 376996 573384 377002 573436
rect 292574 573316 292580 573368
rect 292632 573356 292638 573368
rect 357158 573356 357164 573368
rect 292632 573328 357164 573356
rect 292632 573316 292638 573328
rect 357158 573316 357164 573328
rect 357216 573316 357222 573368
rect 306374 571956 306380 572008
rect 306432 571996 306438 572008
rect 389266 571996 389272 572008
rect 306432 571968 389272 571996
rect 306432 571956 306438 571968
rect 389266 571956 389272 571968
rect 389324 571956 389330 572008
rect 283006 570664 283012 570716
rect 283064 570704 283070 570716
rect 350074 570704 350080 570716
rect 283064 570676 350080 570704
rect 283064 570664 283070 570676
rect 350074 570664 350080 570676
rect 350132 570664 350138 570716
rect 304718 570596 304724 570648
rect 304776 570636 304782 570648
rect 394878 570636 394884 570648
rect 304776 570608 394884 570636
rect 304776 570596 304782 570608
rect 394878 570596 394884 570608
rect 394936 570596 394942 570648
rect 253934 569984 253940 570036
rect 253992 570024 253998 570036
rect 256050 570024 256056 570036
rect 253992 569996 256056 570024
rect 253992 569984 253998 569996
rect 256050 569984 256056 569996
rect 256108 569984 256114 570036
rect 314746 569236 314752 569288
rect 314804 569276 314810 569288
rect 337470 569276 337476 569288
rect 314804 569248 337476 569276
rect 314804 569236 314810 569248
rect 337470 569236 337476 569248
rect 337528 569236 337534 569288
rect 253382 569168 253388 569220
rect 253440 569208 253446 569220
rect 512086 569208 512092 569220
rect 253440 569180 512092 569208
rect 253440 569168 253446 569180
rect 512086 569168 512092 569180
rect 512144 569168 512150 569220
rect 388622 568556 388628 568608
rect 388680 568596 388686 568608
rect 393406 568596 393412 568608
rect 388680 568568 393412 568596
rect 388680 568556 388686 568568
rect 393406 568556 393412 568568
rect 393464 568556 393470 568608
rect 355870 567808 355876 567860
rect 355928 567848 355934 567860
rect 367094 567848 367100 567860
rect 355928 567820 367100 567848
rect 355928 567808 355934 567820
rect 367094 567808 367100 567820
rect 367152 567808 367158 567860
rect 358170 566516 358176 566568
rect 358228 566556 358234 566568
rect 394786 566556 394792 566568
rect 358228 566528 394792 566556
rect 358228 566516 358234 566528
rect 394786 566516 394792 566528
rect 394844 566516 394850 566568
rect 304994 566448 305000 566500
rect 305052 566488 305058 566500
rect 365898 566488 365904 566500
rect 305052 566460 365904 566488
rect 305052 566448 305058 566460
rect 365898 566448 365904 566460
rect 365956 566448 365962 566500
rect 385126 565496 385132 565548
rect 385184 565536 385190 565548
rect 391934 565536 391940 565548
rect 385184 565508 391940 565536
rect 385184 565496 385190 565508
rect 391934 565496 391940 565508
rect 391992 565496 391998 565548
rect 296714 565156 296720 565208
rect 296772 565196 296778 565208
rect 367370 565196 367376 565208
rect 296772 565168 367376 565196
rect 296772 565156 296778 565168
rect 367370 565156 367376 565168
rect 367428 565156 367434 565208
rect 253290 565088 253296 565140
rect 253348 565128 253354 565140
rect 381078 565128 381084 565140
rect 253348 565100 381084 565128
rect 253348 565088 253354 565100
rect 381078 565088 381084 565100
rect 381136 565088 381142 565140
rect 300118 563728 300124 563780
rect 300176 563768 300182 563780
rect 367186 563768 367192 563780
rect 300176 563740 367192 563768
rect 300176 563728 300182 563740
rect 367186 563728 367192 563740
rect 367244 563728 367250 563780
rect 254578 563660 254584 563712
rect 254636 563700 254642 563712
rect 320174 563700 320180 563712
rect 254636 563672 320180 563700
rect 254636 563660 254642 563672
rect 320174 563660 320180 563672
rect 320232 563660 320238 563712
rect 359090 563660 359096 563712
rect 359148 563700 359154 563712
rect 380986 563700 380992 563712
rect 359148 563672 380992 563700
rect 359148 563660 359154 563672
rect 380986 563660 380992 563672
rect 381044 563660 381050 563712
rect 358078 562436 358084 562488
rect 358136 562476 358142 562488
rect 390554 562476 390560 562488
rect 358136 562448 390560 562476
rect 358136 562436 358142 562448
rect 390554 562436 390560 562448
rect 390612 562436 390618 562488
rect 300762 562368 300768 562420
rect 300820 562408 300826 562420
rect 363046 562408 363052 562420
rect 300820 562380 363052 562408
rect 300820 562368 300826 562380
rect 363046 562368 363052 562380
rect 363104 562368 363110 562420
rect 372798 562368 372804 562420
rect 372856 562408 372862 562420
rect 383838 562408 383844 562420
rect 372856 562380 383844 562408
rect 372856 562368 372862 562380
rect 383838 562368 383844 562380
rect 383896 562368 383902 562420
rect 291838 562300 291844 562352
rect 291896 562340 291902 562352
rect 375374 562340 375380 562352
rect 291896 562312 375380 562340
rect 291896 562300 291902 562312
rect 375374 562300 375380 562312
rect 375432 562300 375438 562352
rect 321094 561076 321100 561128
rect 321152 561116 321158 561128
rect 402146 561116 402152 561128
rect 321152 561088 402152 561116
rect 321152 561076 321158 561088
rect 402146 561076 402152 561088
rect 402204 561076 402210 561128
rect 304810 561008 304816 561060
rect 304868 561048 304874 561060
rect 399938 561048 399944 561060
rect 304868 561020 399944 561048
rect 304868 561008 304874 561020
rect 399938 561008 399944 561020
rect 399996 561008 400002 561060
rect 289078 560940 289084 560992
rect 289136 560980 289142 560992
rect 386690 560980 386696 560992
rect 289136 560952 386696 560980
rect 289136 560940 289142 560952
rect 386690 560940 386696 560952
rect 386748 560940 386754 560992
rect 362954 559648 362960 559700
rect 363012 559688 363018 559700
rect 374086 559688 374092 559700
rect 363012 559660 374092 559688
rect 363012 559648 363018 559660
rect 374086 559648 374092 559660
rect 374144 559648 374150 559700
rect 358262 559580 358268 559632
rect 358320 559620 358326 559632
rect 386506 559620 386512 559632
rect 358320 559592 386512 559620
rect 358320 559580 358326 559592
rect 386506 559580 386512 559592
rect 386564 559580 386570 559632
rect 265618 559512 265624 559564
rect 265676 559552 265682 559564
rect 483106 559552 483112 559564
rect 265676 559524 483112 559552
rect 265676 559512 265682 559524
rect 483106 559512 483112 559524
rect 483164 559512 483170 559564
rect 365806 558832 365812 558884
rect 365864 558872 365870 558884
rect 371602 558872 371608 558884
rect 365864 558844 371608 558872
rect 365864 558832 365870 558844
rect 371602 558832 371608 558844
rect 371660 558832 371666 558884
rect 358998 558288 359004 558340
rect 359056 558328 359062 558340
rect 381170 558328 381176 558340
rect 359056 558300 381176 558328
rect 359056 558288 359062 558300
rect 381170 558288 381176 558300
rect 381228 558288 381234 558340
rect 362586 558220 362592 558272
rect 362644 558260 362650 558272
rect 373994 558260 374000 558272
rect 362644 558232 374000 558260
rect 362644 558220 362650 558232
rect 373994 558220 374000 558232
rect 374052 558220 374058 558272
rect 376846 558220 376852 558272
rect 376904 558260 376910 558272
rect 538858 558260 538864 558272
rect 376904 558232 538864 558260
rect 376904 558220 376910 558232
rect 538858 558220 538864 558232
rect 538916 558220 538922 558272
rect 264330 558152 264336 558204
rect 264388 558192 264394 558204
rect 512270 558192 512276 558204
rect 264388 558164 512276 558192
rect 264388 558152 264394 558164
rect 512270 558152 512276 558164
rect 512328 558152 512334 558204
rect 254578 557540 254584 557592
rect 254636 557580 254642 557592
rect 265618 557580 265624 557592
rect 254636 557552 265624 557580
rect 254636 557540 254642 557552
rect 265618 557540 265624 557552
rect 265676 557540 265682 557592
rect 372706 557540 372712 557592
rect 372764 557580 372770 557592
rect 404354 557580 404360 557592
rect 372764 557552 404360 557580
rect 372764 557540 372770 557552
rect 404354 557540 404360 557552
rect 404412 557540 404418 557592
rect 355226 556996 355232 557048
rect 355284 557036 355290 557048
rect 372706 557036 372712 557048
rect 355284 557008 372712 557036
rect 355284 556996 355290 557008
rect 372706 556996 372712 557008
rect 372764 556996 372770 557048
rect 359366 556860 359372 556912
rect 359424 556900 359430 556912
rect 379606 556900 379612 556912
rect 359424 556872 379612 556900
rect 359424 556860 359430 556872
rect 379606 556860 379612 556872
rect 379664 556860 379670 556912
rect 358354 556792 358360 556844
rect 358412 556832 358418 556844
rect 396074 556832 396080 556844
rect 358412 556804 396080 556832
rect 358412 556792 358418 556804
rect 396074 556792 396080 556804
rect 396132 556792 396138 556844
rect 359274 555500 359280 555552
rect 359332 555540 359338 555552
rect 385034 555540 385040 555552
rect 359332 555512 385040 555540
rect 359332 555500 359338 555512
rect 385034 555500 385040 555512
rect 385092 555500 385098 555552
rect 253198 555432 253204 555484
rect 253256 555472 253262 555484
rect 511994 555472 512000 555484
rect 253256 555444 512000 555472
rect 253256 555432 253262 555444
rect 511994 555432 512000 555444
rect 512052 555432 512058 555484
rect 369854 554752 369860 554804
rect 369912 554792 369918 554804
rect 403066 554792 403072 554804
rect 369912 554764 403072 554792
rect 369912 554752 369918 554764
rect 403066 554752 403072 554764
rect 403124 554752 403130 554804
rect 355686 554072 355692 554124
rect 355744 554112 355750 554124
rect 369854 554112 369860 554124
rect 355744 554084 369860 554112
rect 355744 554072 355750 554084
rect 369854 554072 369860 554084
rect 369912 554072 369918 554124
rect 295518 554004 295524 554056
rect 295576 554044 295582 554056
rect 404814 554044 404820 554056
rect 295576 554016 404820 554044
rect 295576 554004 295582 554016
rect 404814 554004 404820 554016
rect 404872 554004 404878 554056
rect 358722 553392 358728 553444
rect 358780 553432 358786 553444
rect 361022 553432 361028 553444
rect 358780 553404 361028 553432
rect 358780 553392 358786 553404
rect 361022 553392 361028 553404
rect 361080 553392 361086 553444
rect 376846 553324 376852 553376
rect 376904 553364 376910 553376
rect 377766 553364 377772 553376
rect 376904 553336 377772 553364
rect 376904 553324 376910 553336
rect 377766 553324 377772 553336
rect 377824 553324 377830 553376
rect 392578 553324 392584 553376
rect 392636 553364 392642 553376
rect 394142 553364 394148 553376
rect 392636 553336 394148 553364
rect 392636 553324 392642 553336
rect 394142 553324 394148 553336
rect 394200 553324 394206 553376
rect 360102 553052 360108 553104
rect 360160 553092 360166 553104
rect 378686 553092 378692 553104
rect 360160 553064 378692 553092
rect 360160 553052 360166 553064
rect 378686 553052 378692 553064
rect 378744 553052 378750 553104
rect 356882 552984 356888 553036
rect 356940 553024 356946 553036
rect 376754 553024 376760 553036
rect 356940 552996 376760 553024
rect 356940 552984 356946 552996
rect 376754 552984 376760 552996
rect 376812 552984 376818 553036
rect 392854 552984 392860 553036
rect 392912 553024 392918 553036
rect 398926 553024 398932 553036
rect 392912 552996 398932 553024
rect 392912 552984 392918 552996
rect 398926 552984 398932 552996
rect 398984 552984 398990 553036
rect 356974 552916 356980 552968
rect 357032 552956 357038 552968
rect 396350 552956 396356 552968
rect 357032 552928 396356 552956
rect 357032 552916 357038 552928
rect 396350 552916 396356 552928
rect 396408 552916 396414 552968
rect 322290 552848 322296 552900
rect 322348 552888 322354 552900
rect 364518 552888 364524 552900
rect 322348 552860 364524 552888
rect 322348 552848 322354 552860
rect 364518 552848 364524 552860
rect 364576 552848 364582 552900
rect 389634 552848 389640 552900
rect 389692 552888 389698 552900
rect 400398 552888 400404 552900
rect 389692 552860 400404 552888
rect 389692 552848 389698 552860
rect 400398 552848 400404 552860
rect 400456 552848 400462 552900
rect 309226 552780 309232 552832
rect 309284 552820 309290 552832
rect 360654 552820 360660 552832
rect 309284 552792 360660 552820
rect 309284 552780 309290 552792
rect 360654 552780 360660 552792
rect 360712 552780 360718 552832
rect 361482 552780 361488 552832
rect 361540 552820 361546 552832
rect 374178 552820 374184 552832
rect 361540 552792 374184 552820
rect 361540 552780 361546 552792
rect 374178 552780 374184 552792
rect 374236 552780 374242 552832
rect 376110 552780 376116 552832
rect 376168 552820 376174 552832
rect 399018 552820 399024 552832
rect 376168 552792 399024 552820
rect 376168 552780 376174 552792
rect 399018 552780 399024 552792
rect 399076 552780 399082 552832
rect 322198 552712 322204 552764
rect 322256 552752 322262 552764
rect 380618 552752 380624 552764
rect 322256 552724 380624 552752
rect 322256 552712 322262 552724
rect 380618 552712 380624 552724
rect 380676 552712 380682 552764
rect 383746 552712 383752 552764
rect 383804 552752 383810 552764
rect 399478 552752 399484 552764
rect 383804 552724 399484 552752
rect 383804 552712 383810 552724
rect 399478 552712 399484 552724
rect 399536 552712 399542 552764
rect 325050 552644 325056 552696
rect 325108 552684 325114 552696
rect 397362 552684 397368 552696
rect 325108 552656 397368 552684
rect 325108 552644 325114 552656
rect 397362 552644 397368 552656
rect 397420 552644 397426 552696
rect 393498 552440 393504 552492
rect 393556 552480 393562 552492
rect 399110 552480 399116 552492
rect 393556 552452 399116 552480
rect 393556 552440 393562 552452
rect 399110 552440 399116 552452
rect 399168 552440 399174 552492
rect 356054 552372 356060 552424
rect 356112 552412 356118 552424
rect 371878 552412 371884 552424
rect 356112 552384 371884 552412
rect 356112 552372 356118 552384
rect 371878 552372 371884 552384
rect 371936 552372 371942 552424
rect 385770 552412 385776 552424
rect 383672 552384 385776 552412
rect 355778 552304 355784 552356
rect 355836 552344 355842 552356
rect 381538 552344 381544 552356
rect 355836 552316 381544 552344
rect 355836 552304 355842 552316
rect 381538 552304 381544 552316
rect 381596 552304 381602 552356
rect 354950 552236 354956 552288
rect 355008 552276 355014 552288
rect 383672 552276 383700 552384
rect 385770 552372 385776 552384
rect 385828 552372 385834 552424
rect 387978 552344 387984 552356
rect 355008 552248 383700 552276
rect 384408 552316 387984 552344
rect 355008 552236 355014 552248
rect 348418 552168 348424 552220
rect 348476 552208 348482 552220
rect 384408 552208 384436 552316
rect 387978 552304 387984 552316
rect 388036 552304 388042 552356
rect 396718 552236 396724 552288
rect 396776 552276 396782 552288
rect 398006 552276 398012 552288
rect 396776 552248 398012 552276
rect 396776 552236 396782 552248
rect 398006 552236 398012 552248
rect 398064 552236 398070 552288
rect 398650 552236 398656 552288
rect 398708 552276 398714 552288
rect 418798 552276 418804 552288
rect 398708 552248 418804 552276
rect 398708 552236 398714 552248
rect 418798 552236 418804 552248
rect 418856 552236 418862 552288
rect 348476 552180 384436 552208
rect 348476 552168 348482 552180
rect 384482 552168 384488 552220
rect 384540 552208 384546 552220
rect 385678 552208 385684 552220
rect 384540 552180 385684 552208
rect 384540 552168 384546 552180
rect 385678 552168 385684 552180
rect 385736 552168 385742 552220
rect 394786 552168 394792 552220
rect 394844 552208 394850 552220
rect 430574 552208 430580 552220
rect 394844 552180 430580 552208
rect 394844 552168 394850 552180
rect 430574 552168 430580 552180
rect 430632 552168 430638 552220
rect 367094 552100 367100 552152
rect 367152 552140 367158 552152
rect 414658 552140 414664 552152
rect 367152 552112 414664 552140
rect 367152 552100 367158 552112
rect 414658 552100 414664 552112
rect 414716 552100 414722 552152
rect 373534 552032 373540 552084
rect 373592 552072 373598 552084
rect 420178 552072 420184 552084
rect 373592 552044 420184 552072
rect 373592 552032 373598 552044
rect 420178 552032 420184 552044
rect 420236 552032 420242 552084
rect 393314 551964 393320 552016
rect 393372 552004 393378 552016
rect 400582 552004 400588 552016
rect 393372 551976 400588 552004
rect 393372 551964 393378 551976
rect 400582 551964 400588 551976
rect 400640 551964 400646 552016
rect 389174 551692 389180 551744
rect 389232 551732 389238 551744
rect 399846 551732 399852 551744
rect 389232 551704 399852 551732
rect 389232 551692 389238 551704
rect 399846 551692 399852 551704
rect 399904 551692 399910 551744
rect 383654 551624 383660 551676
rect 383712 551664 383718 551676
rect 400030 551664 400036 551676
rect 383712 551636 400036 551664
rect 383712 551624 383718 551636
rect 400030 551624 400036 551636
rect 400088 551624 400094 551676
rect 363230 551556 363236 551608
rect 363288 551596 363294 551608
rect 400398 551596 400404 551608
rect 363288 551568 400404 551596
rect 363288 551556 363294 551568
rect 400398 551556 400404 551568
rect 400456 551556 400462 551608
rect 360102 551488 360108 551540
rect 360160 551528 360166 551540
rect 444374 551528 444380 551540
rect 360160 551500 444380 551528
rect 360160 551488 360166 551500
rect 444374 551488 444380 551500
rect 444432 551488 444438 551540
rect 295334 551420 295340 551472
rect 295392 551460 295398 551472
rect 402974 551460 402980 551472
rect 295392 551432 402980 551460
rect 295392 551420 295398 551432
rect 402974 551420 402980 551432
rect 403032 551420 403038 551472
rect 295426 551352 295432 551404
rect 295484 551392 295490 551404
rect 404446 551392 404452 551404
rect 295484 551364 404452 551392
rect 295484 551352 295490 551364
rect 404446 551352 404452 551364
rect 404504 551352 404510 551404
rect 254394 551284 254400 551336
rect 254452 551324 254458 551336
rect 268378 551324 268384 551336
rect 254452 551296 268384 551324
rect 254452 551284 254458 551296
rect 268378 551284 268384 551296
rect 268436 551284 268442 551336
rect 291194 551284 291200 551336
rect 291252 551324 291258 551336
rect 403434 551324 403440 551336
rect 291252 551296 403440 551324
rect 291252 551284 291258 551296
rect 403434 551284 403440 551296
rect 403492 551284 403498 551336
rect 382274 551216 382280 551268
rect 382332 551256 382338 551268
rect 382918 551256 382924 551268
rect 382332 551228 382924 551256
rect 382332 551216 382338 551228
rect 382918 551216 382924 551228
rect 382976 551216 382982 551268
rect 354214 551080 354220 551132
rect 354272 551120 354278 551132
rect 388622 551120 388628 551132
rect 354272 551092 388628 551120
rect 354272 551080 354278 551092
rect 388622 551080 388628 551092
rect 388680 551120 388686 551132
rect 388990 551120 388996 551132
rect 388680 551092 388996 551120
rect 388680 551080 388686 551092
rect 388990 551080 388996 551092
rect 389048 551080 389054 551132
rect 377398 551012 377404 551064
rect 377456 551052 377462 551064
rect 377950 551052 377956 551064
rect 377456 551024 377956 551052
rect 377456 551012 377462 551024
rect 377950 551012 377956 551024
rect 378008 551052 378014 551064
rect 403526 551052 403532 551064
rect 378008 551024 403532 551052
rect 378008 551012 378014 551024
rect 403526 551012 403532 551024
rect 403584 551012 403590 551064
rect 351454 550944 351460 550996
rect 351512 550984 351518 550996
rect 384482 550984 384488 550996
rect 351512 550956 384488 550984
rect 351512 550944 351518 550956
rect 384482 550944 384488 550956
rect 384540 550944 384546 550996
rect 355502 550876 355508 550928
rect 355560 550916 355566 550928
rect 397454 550916 397460 550928
rect 355560 550888 397460 550916
rect 355560 550876 355566 550888
rect 397454 550876 397460 550888
rect 397512 550876 397518 550928
rect 355594 550808 355600 550860
rect 355652 550848 355658 550860
rect 404538 550848 404544 550860
rect 355652 550820 404544 550848
rect 355652 550808 355658 550820
rect 404538 550808 404544 550820
rect 404596 550808 404602 550860
rect 345842 550740 345848 550792
rect 345900 550780 345906 550792
rect 364426 550780 364432 550792
rect 345900 550752 364432 550780
rect 345900 550740 345906 550752
rect 364426 550740 364432 550752
rect 364484 550780 364490 550792
rect 396074 550780 396080 550792
rect 364484 550752 396080 550780
rect 364484 550740 364490 550752
rect 396074 550740 396080 550752
rect 396132 550740 396138 550792
rect 333330 550672 333336 550724
rect 333388 550712 333394 550724
rect 333882 550712 333888 550724
rect 333388 550684 333888 550712
rect 333388 550672 333394 550684
rect 333882 550672 333888 550684
rect 333940 550712 333946 550724
rect 404906 550712 404912 550724
rect 333940 550684 404912 550712
rect 333940 550672 333946 550684
rect 404906 550672 404912 550684
rect 404964 550672 404970 550724
rect 356974 550604 356980 550656
rect 357032 550644 357038 550656
rect 361114 550644 361120 550656
rect 357032 550616 361120 550644
rect 357032 550604 357038 550616
rect 361114 550604 361120 550616
rect 361172 550604 361178 550656
rect 391198 550604 391204 550656
rect 391256 550644 391262 550656
rect 475838 550644 475844 550656
rect 391256 550616 475844 550644
rect 391256 550604 391262 550616
rect 475838 550604 475844 550616
rect 475896 550604 475902 550656
rect 399754 550536 399760 550588
rect 399812 550576 399818 550588
rect 402054 550576 402060 550588
rect 399812 550548 402060 550576
rect 399812 550536 399818 550548
rect 402054 550536 402060 550548
rect 402112 550536 402118 550588
rect 397546 550468 397552 550520
rect 397604 550508 397610 550520
rect 400674 550508 400680 550520
rect 397604 550480 400680 550508
rect 397604 550468 397610 550480
rect 400674 550468 400680 550480
rect 400732 550468 400738 550520
rect 386598 550264 386604 550316
rect 386656 550304 386662 550316
rect 387058 550304 387064 550316
rect 386656 550276 387064 550304
rect 386656 550264 386662 550276
rect 387058 550264 387064 550276
rect 387116 550264 387122 550316
rect 356882 550128 356888 550180
rect 356940 550168 356946 550180
rect 362954 550168 362960 550180
rect 356940 550140 362960 550168
rect 356940 550128 356946 550140
rect 362954 550128 362960 550140
rect 363012 550128 363018 550180
rect 355134 550060 355140 550112
rect 355192 550100 355198 550112
rect 362586 550100 362592 550112
rect 355192 550072 362592 550100
rect 355192 550060 355198 550072
rect 362586 550060 362592 550072
rect 362644 550060 362650 550112
rect 352466 549992 352472 550044
rect 352524 550032 352530 550044
rect 377950 550032 377956 550044
rect 352524 550004 377956 550032
rect 352524 549992 352530 550004
rect 377950 549992 377956 550004
rect 378008 549992 378014 550044
rect 394694 550032 394700 550044
rect 379486 550004 394700 550032
rect 355042 549924 355048 549976
rect 355100 549964 355106 549976
rect 379486 549964 379514 550004
rect 394694 549992 394700 550004
rect 394752 550032 394758 550044
rect 400766 550032 400772 550044
rect 394752 550004 400772 550032
rect 394752 549992 394758 550004
rect 400766 549992 400772 550004
rect 400824 549992 400830 550044
rect 355100 549936 379514 549964
rect 355100 549924 355106 549936
rect 322198 549856 322204 549908
rect 322256 549896 322262 549908
rect 397638 549896 397644 549908
rect 322256 549868 397644 549896
rect 322256 549856 322262 549868
rect 397638 549856 397644 549868
rect 397696 549896 397702 549908
rect 402422 549896 402428 549908
rect 397696 549868 402428 549896
rect 397696 549856 397702 549868
rect 402422 549856 402428 549868
rect 402480 549856 402486 549908
rect 364886 549828 364892 549840
rect 364306 549800 364892 549828
rect 364306 549556 364334 549800
rect 364886 549788 364892 549800
rect 364944 549788 364950 549840
rect 371326 549788 371332 549840
rect 371384 549788 371390 549840
rect 383654 549828 383660 549840
rect 373966 549800 383660 549828
rect 350506 549528 364334 549556
rect 345750 549380 345756 549432
rect 345808 549420 345814 549432
rect 350506 549420 350534 549528
rect 353202 549448 353208 549500
rect 353260 549488 353266 549500
rect 371344 549488 371372 549788
rect 353260 549460 371372 549488
rect 353260 549448 353266 549460
rect 345808 549392 350534 549420
rect 345808 549380 345814 549392
rect 326982 549312 326988 549364
rect 327040 549352 327046 549364
rect 355134 549352 355140 549364
rect 327040 549324 355140 549352
rect 327040 549312 327046 549324
rect 355134 549312 355140 549324
rect 355192 549312 355198 549364
rect 325050 549244 325056 549296
rect 325108 549284 325114 549296
rect 373966 549284 373994 549800
rect 383654 549788 383660 549800
rect 383712 549788 383718 549840
rect 325108 549256 373994 549284
rect 325108 549244 325114 549256
rect 322290 548564 322296 548616
rect 322348 548604 322354 548616
rect 356054 548604 356060 548616
rect 322348 548576 356060 548604
rect 322348 548564 322354 548576
rect 356054 548564 356060 548576
rect 356112 548564 356118 548616
rect 304902 548496 304908 548548
rect 304960 548536 304966 548548
rect 341518 548536 341524 548548
rect 304960 548508 341524 548536
rect 304960 548496 304966 548508
rect 341518 548496 341524 548508
rect 341576 548496 341582 548548
rect 281534 547816 281540 547868
rect 281592 547856 281598 547868
rect 357434 547856 357440 547868
rect 281592 547828 357440 547856
rect 281592 547816 281598 547828
rect 357434 547816 357440 547828
rect 357492 547816 357498 547868
rect 316678 546388 316684 546440
rect 316736 546428 316742 546440
rect 357434 546428 357440 546440
rect 316736 546400 357440 546428
rect 316736 546388 316742 546400
rect 357434 546388 357440 546400
rect 357492 546388 357498 546440
rect 279510 545844 279516 545896
rect 279568 545884 279574 545896
rect 313642 545884 313648 545896
rect 279568 545856 313648 545884
rect 279568 545844 279574 545856
rect 313642 545844 313648 545856
rect 313700 545844 313706 545896
rect 279602 545708 279608 545760
rect 279660 545748 279666 545760
rect 312906 545748 312912 545760
rect 279660 545720 312912 545748
rect 279660 545708 279666 545720
rect 312906 545708 312912 545720
rect 312964 545708 312970 545760
rect 313274 545708 313280 545760
rect 313332 545748 313338 545760
rect 349982 545748 349988 545760
rect 313332 545720 349988 545748
rect 313332 545708 313338 545720
rect 349982 545708 349988 545720
rect 350040 545708 350046 545760
rect 307662 545028 307668 545080
rect 307720 545068 307726 545080
rect 357434 545068 357440 545080
rect 307720 545040 357440 545068
rect 307720 545028 307726 545040
rect 357434 545028 357440 545040
rect 357492 545028 357498 545080
rect 278958 543600 278964 543652
rect 279016 543640 279022 543652
rect 297450 543640 297456 543652
rect 279016 543612 297456 543640
rect 279016 543600 279022 543612
rect 297450 543600 297456 543612
rect 297508 543600 297514 543652
rect 279234 543532 279240 543584
rect 279292 543572 279298 543584
rect 300394 543572 300400 543584
rect 279292 543544 300400 543572
rect 279292 543532 279298 543544
rect 300394 543532 300400 543544
rect 300452 543532 300458 543584
rect 279970 543464 279976 543516
rect 280028 543504 280034 543516
rect 301130 543504 301136 543516
rect 280028 543476 301136 543504
rect 280028 543464 280034 543476
rect 301130 543464 301136 543476
rect 301188 543464 301194 543516
rect 280062 543396 280068 543448
rect 280120 543436 280126 543448
rect 302602 543436 302608 543448
rect 280120 543408 302608 543436
rect 280120 543396 280126 543408
rect 302602 543396 302608 543408
rect 302660 543396 302666 543448
rect 401594 543396 401600 543448
rect 401652 543436 401658 543448
rect 404538 543436 404544 543448
rect 401652 543408 404544 543436
rect 401652 543396 401658 543408
rect 404538 543396 404544 543408
rect 404596 543396 404602 543448
rect 279418 543328 279424 543380
rect 279476 543368 279482 543380
rect 303798 543368 303804 543380
rect 279476 543340 303804 543368
rect 279476 543328 279482 543340
rect 303798 543328 303804 543340
rect 303856 543328 303862 543380
rect 279326 543260 279332 543312
rect 279384 543300 279390 543312
rect 305546 543300 305552 543312
rect 279384 543272 305552 543300
rect 279384 543260 279390 543272
rect 305546 543260 305552 543272
rect 305604 543260 305610 543312
rect 279142 543192 279148 543244
rect 279200 543232 279206 543244
rect 316034 543232 316040 543244
rect 279200 543204 316040 543232
rect 279200 543192 279206 543204
rect 316034 543192 316040 543204
rect 316092 543192 316098 543244
rect 279050 543124 279056 543176
rect 279108 543164 279114 543176
rect 315114 543164 315120 543176
rect 279108 543136 315120 543164
rect 279108 543124 279114 543136
rect 315114 543124 315120 543136
rect 315172 543124 315178 543176
rect 278130 543056 278136 543108
rect 278188 543096 278194 543108
rect 316586 543096 316592 543108
rect 278188 543068 316592 543096
rect 278188 543056 278194 543068
rect 316586 543056 316592 543068
rect 316644 543056 316650 543108
rect 257430 542988 257436 543040
rect 257488 543028 257494 543040
rect 314838 543028 314844 543040
rect 257488 543000 314844 543028
rect 257488 542988 257494 543000
rect 314838 542988 314844 543000
rect 314896 542988 314902 543040
rect 323670 542988 323676 543040
rect 323728 543028 323734 543040
rect 357526 543028 357532 543040
rect 323728 543000 357532 543028
rect 323728 542988 323734 543000
rect 357526 542988 357532 543000
rect 357584 542988 357590 543040
rect 279694 542580 279700 542632
rect 279752 542620 279758 542632
rect 294506 542620 294512 542632
rect 279752 542592 294512 542620
rect 279752 542580 279758 542592
rect 294506 542580 294512 542592
rect 294564 542580 294570 542632
rect 279602 542512 279608 542564
rect 279660 542552 279666 542564
rect 293954 542552 293960 542564
rect 279660 542524 293960 542552
rect 279660 542512 279666 542524
rect 293954 542512 293960 542524
rect 294012 542512 294018 542564
rect 279878 542444 279884 542496
rect 279936 542484 279942 542496
rect 295334 542484 295340 542496
rect 279936 542456 295340 542484
rect 279936 542444 279942 542456
rect 295334 542444 295340 542456
rect 295392 542444 295398 542496
rect 279510 542376 279516 542428
rect 279568 542416 279574 542428
rect 295978 542416 295984 542428
rect 279568 542388 295984 542416
rect 279568 542376 279574 542388
rect 295978 542376 295984 542388
rect 296036 542376 296042 542428
rect 306282 541696 306288 541748
rect 306340 541736 306346 541748
rect 340230 541736 340236 541748
rect 306340 541708 340236 541736
rect 306340 541696 306346 541708
rect 340230 541696 340236 541708
rect 340288 541696 340294 541748
rect 254670 541628 254676 541680
rect 254728 541668 254734 541680
rect 266998 541668 267004 541680
rect 254728 541640 267004 541668
rect 254728 541628 254734 541640
rect 266998 541628 267004 541640
rect 267056 541628 267062 541680
rect 309134 541628 309140 541680
rect 309192 541668 309198 541680
rect 354122 541668 354128 541680
rect 309192 541640 354128 541668
rect 309192 541628 309198 541640
rect 354122 541628 354128 541640
rect 354180 541628 354186 541680
rect 254578 541152 254584 541204
rect 254636 541192 254642 541204
rect 260190 541192 260196 541204
rect 254636 541164 260196 541192
rect 254636 541152 254642 541164
rect 260190 541152 260196 541164
rect 260248 541152 260254 541204
rect 401594 540948 401600 541000
rect 401652 540988 401658 541000
rect 437474 540988 437480 541000
rect 401652 540960 437480 540988
rect 401652 540948 401658 540960
rect 437474 540948 437480 540960
rect 437532 540948 437538 541000
rect 317414 540200 317420 540252
rect 317472 540240 317478 540252
rect 330478 540240 330484 540252
rect 317472 540212 330484 540240
rect 317472 540200 317478 540212
rect 330478 540200 330484 540212
rect 330536 540200 330542 540252
rect 278314 539656 278320 539708
rect 278372 539696 278378 539708
rect 283466 539696 283472 539708
rect 278372 539668 283472 539696
rect 278372 539656 278378 539668
rect 283466 539656 283472 539668
rect 283524 539656 283530 539708
rect 276658 539588 276664 539640
rect 276716 539628 276722 539640
rect 286410 539628 286416 539640
rect 276716 539600 286416 539628
rect 276716 539588 276722 539600
rect 286410 539588 286416 539600
rect 286468 539588 286474 539640
rect 280798 539520 280804 539572
rect 280856 539560 280862 539572
rect 284202 539560 284208 539572
rect 280856 539532 284208 539560
rect 280856 539520 280862 539532
rect 284202 539520 284208 539532
rect 284260 539520 284266 539572
rect 330478 539520 330484 539572
rect 330536 539560 330542 539572
rect 357434 539560 357440 539572
rect 330536 539532 357440 539560
rect 330536 539520 330542 539532
rect 357434 539520 357440 539532
rect 357492 539520 357498 539572
rect 281166 539452 281172 539504
rect 281224 539492 281230 539504
rect 284938 539492 284944 539504
rect 281224 539464 284944 539492
rect 281224 539452 281230 539464
rect 284938 539452 284944 539464
rect 284996 539452 285002 539504
rect 320174 537480 320180 537532
rect 320232 537520 320238 537532
rect 325602 537520 325608 537532
rect 320232 537492 325608 537520
rect 320232 537480 320238 537492
rect 325602 537480 325608 537492
rect 325660 537520 325666 537532
rect 329098 537520 329104 537532
rect 325660 537492 329104 537520
rect 325660 537480 325666 537492
rect 329098 537480 329104 537492
rect 329156 537480 329162 537532
rect 340874 536800 340880 536852
rect 340932 536840 340938 536852
rect 358354 536840 358360 536852
rect 340932 536812 358360 536840
rect 340932 536800 340938 536812
rect 358354 536800 358360 536812
rect 358412 536800 358418 536852
rect 485498 536800 485504 536852
rect 485556 536840 485562 536852
rect 579890 536840 579896 536852
rect 485556 536812 579896 536840
rect 485556 536800 485562 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 349890 536732 349896 536784
rect 349948 536772 349954 536784
rect 357434 536772 357440 536784
rect 349948 536744 357440 536772
rect 349948 536732 349954 536744
rect 357434 536732 357440 536744
rect 357492 536732 357498 536784
rect 355410 536664 355416 536716
rect 355468 536704 355474 536716
rect 357894 536704 357900 536716
rect 355468 536676 357900 536704
rect 355468 536664 355474 536676
rect 357894 536664 357900 536676
rect 357952 536664 357958 536716
rect 401594 536188 401600 536240
rect 401652 536228 401658 536240
rect 403342 536228 403348 536240
rect 401652 536200 403348 536228
rect 401652 536188 401658 536200
rect 403342 536188 403348 536200
rect 403400 536188 403406 536240
rect 322382 536052 322388 536104
rect 322440 536092 322446 536104
rect 340874 536092 340880 536104
rect 322440 536064 340880 536092
rect 322440 536052 322446 536064
rect 340874 536052 340880 536064
rect 340932 536052 340938 536104
rect 477494 536052 477500 536104
rect 477552 536092 477558 536104
rect 502886 536092 502892 536104
rect 477552 536064 502892 536092
rect 477552 536052 477558 536064
rect 502886 536052 502892 536064
rect 502944 536052 502950 536104
rect 338850 535372 338856 535424
rect 338908 535412 338914 535424
rect 357434 535412 357440 535424
rect 338908 535384 357440 535412
rect 338908 535372 338914 535384
rect 357434 535372 357440 535384
rect 357492 535372 357498 535424
rect 350074 535304 350080 535356
rect 350132 535344 350138 535356
rect 357526 535344 357532 535356
rect 350132 535316 357532 535344
rect 350132 535304 350138 535316
rect 357526 535304 357532 535316
rect 357584 535304 357590 535356
rect 353110 535236 353116 535288
rect 353168 535276 353174 535288
rect 357434 535276 357440 535288
rect 353168 535248 357440 535276
rect 353168 535236 353174 535248
rect 357434 535236 357440 535248
rect 357492 535236 357498 535288
rect 322474 534692 322480 534744
rect 322532 534732 322538 534744
rect 330478 534732 330484 534744
rect 322532 534704 330484 534732
rect 322532 534692 322538 534704
rect 330478 534692 330484 534704
rect 330536 534692 330542 534744
rect 254670 534080 254676 534132
rect 254728 534120 254734 534132
rect 278130 534120 278136 534132
rect 254728 534092 278136 534120
rect 254728 534080 254734 534092
rect 278130 534080 278136 534092
rect 278188 534080 278194 534132
rect 322474 534080 322480 534132
rect 322532 534120 322538 534132
rect 359734 534120 359740 534132
rect 322532 534092 359740 534120
rect 322532 534080 322538 534092
rect 359734 534080 359740 534092
rect 359792 534080 359798 534132
rect 401870 533740 401876 533792
rect 401928 533780 401934 533792
rect 404354 533780 404360 533792
rect 401928 533752 404360 533780
rect 401928 533740 401934 533752
rect 404354 533740 404360 533752
rect 404412 533740 404418 533792
rect 358170 533468 358176 533520
rect 358228 533468 358234 533520
rect 322842 533400 322848 533452
rect 322900 533440 322906 533452
rect 340138 533440 340144 533452
rect 322900 533412 340144 533440
rect 322900 533400 322906 533412
rect 340138 533400 340144 533412
rect 340196 533400 340202 533452
rect 328362 533332 328368 533384
rect 328420 533372 328426 533384
rect 357710 533372 357716 533384
rect 328420 533344 357716 533372
rect 328420 533332 328426 533344
rect 357710 533332 357716 533344
rect 357768 533372 357774 533384
rect 358188 533372 358216 533468
rect 357768 533344 358216 533372
rect 357768 533332 357774 533344
rect 481542 533332 481548 533384
rect 481600 533372 481606 533384
rect 526438 533372 526444 533384
rect 481600 533344 526444 533372
rect 481600 533332 481606 533344
rect 526438 533332 526444 533344
rect 526496 533332 526502 533384
rect 323762 532720 323768 532772
rect 323820 532760 323826 532772
rect 350534 532760 350540 532772
rect 323820 532732 350540 532760
rect 323820 532720 323826 532732
rect 350534 532720 350540 532732
rect 350592 532720 350598 532772
rect 321646 532652 321652 532704
rect 321704 532692 321710 532704
rect 355134 532692 355140 532704
rect 321704 532664 355140 532692
rect 321704 532652 321710 532664
rect 355134 532652 355140 532664
rect 355192 532652 355198 532704
rect 327810 532584 327816 532636
rect 327868 532624 327874 532636
rect 357434 532624 357440 532636
rect 327868 532596 357440 532624
rect 327868 532584 327874 532596
rect 357434 532584 357440 532596
rect 357492 532584 357498 532636
rect 335998 532516 336004 532568
rect 336056 532556 336062 532568
rect 357526 532556 357532 532568
rect 336056 532528 357532 532556
rect 336056 532516 336062 532528
rect 357526 532516 357532 532528
rect 357584 532516 357590 532568
rect 350534 532448 350540 532500
rect 350592 532488 350598 532500
rect 351178 532488 351184 532500
rect 350592 532460 351184 532488
rect 350592 532448 350598 532460
rect 351178 532448 351184 532460
rect 351236 532488 351242 532500
rect 355226 532488 355232 532500
rect 351236 532460 355232 532488
rect 351236 532448 351242 532460
rect 355226 532448 355232 532460
rect 355284 532448 355290 532500
rect 475470 531972 475476 532024
rect 475528 532012 475534 532024
rect 492674 532012 492680 532024
rect 475528 531984 492680 532012
rect 475528 531972 475534 531984
rect 492674 531972 492680 531984
rect 492732 531972 492738 532024
rect 494422 531972 494428 532024
rect 494480 532012 494486 532024
rect 582374 532012 582380 532024
rect 494480 531984 582380 532012
rect 494480 531972 494486 531984
rect 582374 531972 582380 531984
rect 582432 531972 582438 532024
rect 401962 531904 401968 531956
rect 402020 531944 402026 531956
rect 404722 531944 404728 531956
rect 402020 531916 404728 531944
rect 402020 531904 402026 531916
rect 404722 531904 404728 531916
rect 404780 531904 404786 531956
rect 434714 531904 434720 531956
rect 434772 531944 434778 531956
rect 505554 531944 505560 531956
rect 434772 531916 505560 531944
rect 434772 531904 434778 531916
rect 505554 531904 505560 531916
rect 505612 531904 505618 531956
rect 416774 531836 416780 531888
rect 416832 531876 416838 531888
rect 497734 531876 497740 531888
rect 416832 531848 497740 531876
rect 416832 531836 416838 531848
rect 497734 531836 497740 531848
rect 497792 531836 497798 531888
rect 438854 531768 438860 531820
rect 438912 531808 438918 531820
rect 496446 531808 496452 531820
rect 438912 531780 496452 531808
rect 438912 531768 438918 531780
rect 496446 531768 496452 531780
rect 496504 531768 496510 531820
rect 475378 531700 475384 531752
rect 475436 531740 475442 531752
rect 506106 531740 506112 531752
rect 475436 531712 506112 531740
rect 475436 531700 475442 531712
rect 506106 531700 506112 531712
rect 506164 531700 506170 531752
rect 507210 531700 507216 531752
rect 507268 531740 507274 531752
rect 549898 531740 549904 531752
rect 507268 531712 549904 531740
rect 507268 531700 507274 531712
rect 549898 531700 549904 531712
rect 549956 531700 549962 531752
rect 476758 531632 476764 531684
rect 476816 531672 476822 531684
rect 508774 531672 508780 531684
rect 476816 531644 508780 531672
rect 476816 531632 476822 531644
rect 508774 531632 508780 531644
rect 508832 531632 508838 531684
rect 463694 531564 463700 531616
rect 463752 531604 463758 531616
rect 495434 531604 495440 531616
rect 463752 531576 495440 531604
rect 463752 531564 463758 531576
rect 495434 531564 495440 531576
rect 495492 531564 495498 531616
rect 499298 531564 499304 531616
rect 499356 531604 499362 531616
rect 527818 531604 527824 531616
rect 499356 531576 527824 531604
rect 499356 531564 499362 531576
rect 527818 531564 527824 531576
rect 527876 531564 527882 531616
rect 448514 531496 448520 531548
rect 448572 531536 448578 531548
rect 487430 531536 487436 531548
rect 448572 531508 487436 531536
rect 448572 531496 448578 531508
rect 487430 531496 487436 531508
rect 487488 531496 487494 531548
rect 504174 531496 504180 531548
rect 504232 531536 504238 531548
rect 534718 531536 534724 531548
rect 504232 531508 534724 531536
rect 504232 531496 504238 531508
rect 534718 531496 534724 531508
rect 534776 531496 534782 531548
rect 476942 531428 476948 531480
rect 477000 531468 477006 531480
rect 488074 531468 488080 531480
rect 477000 531440 488080 531468
rect 477000 531428 477006 531440
rect 488074 531428 488080 531440
rect 488132 531428 488138 531480
rect 508682 531428 508688 531480
rect 508740 531468 508746 531480
rect 538858 531468 538864 531480
rect 508740 531440 538864 531468
rect 508740 531428 508746 531440
rect 538858 531428 538864 531440
rect 538916 531428 538922 531480
rect 473354 531360 473360 531412
rect 473412 531400 473418 531412
rect 486786 531400 486792 531412
rect 473412 531372 486792 531400
rect 473412 531360 473418 531372
rect 486786 531360 486792 531372
rect 486844 531360 486850 531412
rect 493870 531360 493876 531412
rect 493928 531400 493934 531412
rect 509878 531400 509884 531412
rect 493928 531372 509884 531400
rect 493928 531360 493934 531372
rect 509878 531360 509884 531372
rect 509936 531360 509942 531412
rect 476850 531292 476856 531344
rect 476908 531332 476914 531344
rect 483566 531332 483572 531344
rect 476908 531304 483572 531332
rect 476908 531292 476914 531304
rect 483566 531292 483572 531304
rect 483624 531292 483630 531344
rect 505462 531292 505468 531344
rect 505520 531332 505526 531344
rect 510614 531332 510620 531344
rect 505520 531304 510620 531332
rect 505520 531292 505526 531304
rect 510614 531292 510620 531304
rect 510672 531292 510678 531344
rect 401962 531224 401968 531276
rect 402020 531264 402026 531276
rect 404446 531264 404452 531276
rect 402020 531236 404452 531264
rect 402020 531224 402026 531236
rect 404446 531224 404452 531236
rect 404504 531224 404510 531276
rect 322474 531156 322480 531208
rect 322532 531196 322538 531208
rect 328362 531196 328368 531208
rect 322532 531168 328368 531196
rect 322532 531156 322538 531168
rect 328362 531156 328368 531168
rect 328420 531156 328426 531208
rect 485038 530544 485044 530596
rect 485096 530584 485102 530596
rect 491938 530584 491944 530596
rect 485096 530556 491944 530584
rect 485096 530544 485102 530556
rect 491938 530544 491944 530556
rect 491996 530544 492002 530596
rect 407114 530476 407120 530528
rect 407172 530516 407178 530528
rect 495802 530516 495808 530528
rect 407172 530488 495808 530516
rect 407172 530476 407178 530488
rect 495802 530476 495808 530488
rect 495860 530476 495866 530528
rect 475562 530408 475568 530460
rect 475620 530448 475626 530460
rect 494514 530448 494520 530460
rect 475620 530420 494520 530448
rect 475620 530408 475626 530420
rect 494514 530408 494520 530420
rect 494572 530408 494578 530460
rect 478874 530340 478880 530392
rect 478932 530380 478938 530392
rect 500310 530380 500316 530392
rect 478932 530352 500316 530380
rect 478932 530340 478938 530352
rect 500310 530340 500316 530352
rect 500368 530340 500374 530392
rect 357710 530272 357716 530324
rect 357768 530312 357774 530324
rect 359458 530312 359464 530324
rect 357768 530284 359464 530312
rect 357768 530272 357774 530284
rect 359458 530272 359464 530284
rect 359516 530272 359522 530324
rect 468478 530272 468484 530324
rect 468536 530312 468542 530324
rect 485038 530312 485044 530324
rect 468536 530284 485044 530312
rect 468536 530272 468542 530284
rect 485038 530272 485044 530284
rect 485096 530272 485102 530324
rect 472618 530204 472624 530256
rect 472676 530244 472682 530256
rect 497090 530244 497096 530256
rect 472676 530216 497096 530244
rect 472676 530204 472682 530216
rect 497090 530204 497096 530216
rect 497148 530204 497154 530256
rect 485820 530136 485826 530188
rect 485878 530176 485884 530188
rect 563054 530176 563060 530188
rect 485878 530148 563060 530176
rect 485878 530136 485884 530148
rect 563054 530136 563060 530148
rect 563112 530136 563118 530188
rect 409874 530068 409880 530120
rect 409932 530108 409938 530120
rect 491616 530108 491622 530120
rect 409932 530080 491622 530108
rect 409932 530068 409938 530080
rect 491616 530068 491622 530080
rect 491674 530068 491680 530120
rect 359826 530040 359832 530052
rect 354646 530012 359832 530040
rect 322382 529932 322388 529984
rect 322440 529972 322446 529984
rect 354646 529972 354674 530012
rect 359826 530000 359832 530012
rect 359884 530000 359890 530052
rect 402882 530000 402888 530052
rect 402940 530040 402946 530052
rect 458174 530040 458180 530052
rect 402940 530012 458180 530040
rect 402940 530000 402946 530012
rect 458174 530000 458180 530012
rect 458232 530000 458238 530052
rect 480990 530000 480996 530052
rect 481048 530040 481054 530052
rect 565814 530040 565820 530052
rect 481048 530012 565820 530040
rect 481048 530000 481054 530012
rect 565814 530000 565820 530012
rect 565872 530000 565878 530052
rect 322440 529944 354674 529972
rect 322440 529932 322446 529944
rect 400858 529932 400864 529984
rect 400916 529972 400922 529984
rect 401870 529972 401876 529984
rect 400916 529944 401876 529972
rect 400916 529932 400922 529944
rect 401870 529932 401876 529944
rect 401928 529932 401934 529984
rect 491202 529932 491208 529984
rect 491260 529972 491266 529984
rect 571978 529972 571984 529984
rect 491260 529944 571984 529972
rect 491260 529932 491266 529944
rect 571978 529932 571984 529944
rect 572036 529932 572042 529984
rect 322474 529864 322480 529916
rect 322532 529904 322538 529916
rect 354214 529904 354220 529916
rect 322532 529876 354220 529904
rect 322532 529864 322538 529876
rect 354214 529864 354220 529876
rect 354272 529864 354278 529916
rect 406378 529864 406384 529916
rect 406436 529904 406442 529916
rect 477494 529904 477500 529916
rect 406436 529876 477500 529904
rect 406436 529864 406442 529876
rect 477494 529864 477500 529876
rect 477552 529864 477558 529916
rect 337470 529796 337476 529848
rect 337528 529836 337534 529848
rect 357434 529836 357440 529848
rect 337528 529808 357440 529836
rect 337528 529796 337534 529808
rect 357434 529796 357440 529808
rect 357492 529796 357498 529848
rect 322842 529184 322848 529236
rect 322900 529224 322906 529236
rect 337562 529224 337568 529236
rect 322900 529196 337568 529224
rect 322900 529184 322906 529196
rect 337562 529184 337568 529196
rect 337620 529184 337626 529236
rect 509786 528844 509792 528896
rect 509844 528884 509850 528896
rect 513374 528884 513380 528896
rect 509844 528856 513380 528884
rect 509844 528844 509850 528856
rect 513374 528844 513380 528856
rect 513432 528844 513438 528896
rect 254210 528572 254216 528624
rect 254268 528612 254274 528624
rect 269850 528612 269856 528624
rect 254268 528584 269856 528612
rect 254268 528572 254274 528584
rect 269850 528572 269856 528584
rect 269908 528572 269914 528624
rect 402882 528572 402888 528624
rect 402940 528612 402946 528624
rect 409138 528612 409144 528624
rect 402940 528584 409144 528612
rect 402940 528572 402946 528584
rect 409138 528572 409144 528584
rect 409196 528572 409202 528624
rect 416038 528572 416044 528624
rect 416096 528612 416102 528624
rect 477494 528612 477500 528624
rect 416096 528584 477500 528612
rect 416096 528572 416102 528584
rect 477494 528572 477500 528584
rect 477552 528572 477558 528624
rect 513282 528572 513288 528624
rect 513340 528612 513346 528624
rect 518158 528612 518164 528624
rect 513340 528584 518164 528612
rect 513340 528572 513346 528584
rect 518158 528572 518164 528584
rect 518216 528572 518222 528624
rect 322474 528504 322480 528556
rect 322532 528544 322538 528556
rect 356974 528544 356980 528556
rect 322532 528516 356980 528544
rect 322532 528504 322538 528516
rect 356974 528504 356980 528516
rect 357032 528504 357038 528556
rect 401962 528300 401968 528352
rect 402020 528340 402026 528352
rect 404630 528340 404636 528352
rect 402020 528312 404636 528340
rect 402020 528300 402026 528312
rect 404630 528300 404636 528312
rect 404688 528300 404694 528352
rect 509878 527824 509884 527876
rect 509936 527864 509942 527876
rect 569954 527864 569960 527876
rect 509936 527836 569960 527864
rect 509936 527824 509942 527836
rect 569954 527824 569960 527836
rect 570012 527824 570018 527876
rect 321554 527212 321560 527264
rect 321612 527252 321618 527264
rect 323670 527252 323676 527264
rect 321612 527224 323676 527252
rect 321612 527212 321618 527224
rect 323670 527212 323676 527224
rect 323728 527212 323734 527264
rect 420914 527144 420920 527196
rect 420972 527184 420978 527196
rect 477494 527184 477500 527196
rect 420972 527156 477500 527184
rect 420972 527144 420978 527156
rect 477494 527144 477500 527156
rect 477552 527144 477558 527196
rect 322474 527076 322480 527128
rect 322532 527116 322538 527128
rect 351454 527116 351460 527128
rect 322532 527088 351460 527116
rect 322532 527076 322538 527088
rect 351454 527076 351460 527088
rect 351512 527076 351518 527128
rect 355318 527076 355324 527128
rect 355376 527116 355382 527128
rect 357894 527116 357900 527128
rect 355376 527088 357900 527116
rect 355376 527076 355382 527088
rect 357894 527076 357900 527088
rect 357952 527076 357958 527128
rect 331858 527008 331864 527060
rect 331916 527048 331922 527060
rect 357434 527048 357440 527060
rect 331916 527020 357440 527048
rect 331916 527008 331922 527020
rect 357434 527008 357440 527020
rect 357492 527008 357498 527060
rect 402238 526736 402244 526788
rect 402296 526776 402302 526788
rect 405090 526776 405096 526788
rect 402296 526748 405096 526776
rect 402296 526736 402302 526748
rect 405090 526736 405096 526748
rect 405148 526736 405154 526788
rect 401778 526396 401784 526448
rect 401836 526436 401842 526448
rect 478874 526436 478880 526448
rect 401836 526408 478880 526436
rect 401836 526396 401842 526408
rect 478874 526396 478880 526408
rect 478932 526396 478938 526448
rect 405090 525784 405096 525836
rect 405148 525824 405154 525836
rect 477494 525824 477500 525836
rect 405148 525796 477500 525824
rect 405148 525784 405154 525796
rect 477494 525784 477500 525796
rect 477552 525784 477558 525836
rect 322474 525716 322480 525768
rect 322532 525756 322538 525768
rect 355042 525756 355048 525768
rect 322532 525728 355048 525756
rect 322532 525716 322538 525728
rect 355042 525716 355048 525728
rect 355100 525716 355106 525768
rect 399662 525716 399668 525768
rect 399720 525756 399726 525768
rect 402422 525756 402428 525768
rect 399720 525728 402428 525756
rect 399720 525716 399726 525728
rect 402422 525716 402428 525728
rect 402480 525716 402486 525768
rect 422938 525716 422944 525768
rect 422996 525756 423002 525768
rect 478690 525756 478696 525768
rect 422996 525728 478696 525756
rect 422996 525716 423002 525728
rect 478690 525716 478696 525728
rect 478748 525716 478754 525768
rect 530578 525716 530584 525768
rect 530636 525756 530642 525768
rect 580166 525756 580172 525768
rect 530636 525728 580172 525756
rect 530636 525716 530642 525728
rect 580166 525716 580172 525728
rect 580224 525716 580230 525768
rect 475746 525580 475752 525632
rect 475804 525620 475810 525632
rect 477954 525620 477960 525632
rect 475804 525592 477960 525620
rect 475804 525580 475810 525592
rect 477954 525580 477960 525592
rect 478012 525580 478018 525632
rect 402238 525308 402244 525360
rect 402296 525348 402302 525360
rect 404906 525348 404912 525360
rect 402296 525320 404912 525348
rect 402296 525308 402302 525320
rect 404906 525308 404912 525320
rect 404964 525308 404970 525360
rect 322750 525036 322756 525088
rect 322808 525076 322814 525088
rect 349890 525076 349896 525088
rect 322808 525048 349896 525076
rect 322808 525036 322814 525048
rect 349890 525036 349896 525048
rect 349948 525036 349954 525088
rect 512638 524424 512644 524476
rect 512696 524464 512702 524476
rect 525058 524464 525064 524476
rect 512696 524436 525064 524464
rect 512696 524424 512702 524436
rect 525058 524424 525064 524436
rect 525116 524424 525122 524476
rect 333238 524356 333244 524408
rect 333296 524396 333302 524408
rect 357434 524396 357440 524408
rect 333296 524368 357440 524396
rect 333296 524356 333302 524368
rect 357434 524356 357440 524368
rect 357492 524356 357498 524408
rect 471330 523200 471336 523252
rect 471388 523240 471394 523252
rect 477494 523240 477500 523252
rect 471388 523212 477500 523240
rect 471388 523200 471394 523212
rect 477494 523200 477500 523212
rect 477552 523200 477558 523252
rect 254026 522996 254032 523048
rect 254084 523036 254090 523048
rect 275370 523036 275376 523048
rect 254084 523008 275376 523036
rect 254084 522996 254090 523008
rect 275370 522996 275376 523008
rect 275428 522996 275434 523048
rect 322474 522996 322480 523048
rect 322532 523036 322538 523048
rect 355870 523036 355876 523048
rect 322532 523008 355876 523036
rect 322532 522996 322538 523008
rect 355870 522996 355876 523008
rect 355928 522996 355934 523048
rect 456794 522996 456800 523048
rect 456852 523036 456858 523048
rect 477494 523036 477500 523048
rect 456852 523008 477500 523036
rect 456852 522996 456858 523008
rect 477494 522996 477500 523008
rect 477552 522996 477558 523048
rect 322014 522928 322020 522980
rect 322072 522968 322078 522980
rect 355778 522968 355784 522980
rect 322072 522940 355784 522968
rect 322072 522928 322078 522940
rect 355778 522928 355784 522940
rect 355836 522928 355842 522980
rect 357618 522928 357624 522980
rect 357676 522968 357682 522980
rect 359642 522968 359648 522980
rect 357676 522940 359648 522968
rect 357676 522928 357682 522940
rect 359642 522928 359648 522940
rect 359700 522928 359706 522980
rect 322474 521636 322480 521688
rect 322532 521676 322538 521688
rect 351454 521676 351460 521688
rect 322532 521648 351460 521676
rect 322532 521636 322538 521648
rect 351454 521636 351460 521648
rect 351512 521636 351518 521688
rect 402882 521636 402888 521688
rect 402940 521676 402946 521688
rect 423674 521676 423680 521688
rect 402940 521648 423680 521676
rect 402940 521636 402946 521648
rect 423674 521636 423680 521648
rect 423732 521636 423738 521688
rect 322014 521568 322020 521620
rect 322072 521608 322078 521620
rect 352466 521608 352472 521620
rect 322072 521580 352472 521608
rect 322072 521568 322078 521580
rect 352466 521568 352472 521580
rect 352524 521568 352530 521620
rect 352466 521024 352472 521076
rect 352524 521064 352530 521076
rect 353294 521064 353300 521076
rect 352524 521036 353300 521064
rect 352524 521024 352530 521036
rect 353294 521024 353300 521036
rect 353352 521024 353358 521076
rect 401594 520956 401600 521008
rect 401652 520996 401658 521008
rect 403526 520996 403532 521008
rect 401652 520968 403532 520996
rect 401652 520956 401658 520968
rect 403526 520956 403532 520968
rect 403584 520956 403590 521008
rect 322474 520276 322480 520328
rect 322532 520316 322538 520328
rect 353110 520316 353116 520328
rect 322532 520288 353116 520316
rect 322532 520276 322538 520288
rect 353110 520276 353116 520288
rect 353168 520276 353174 520328
rect 450538 520276 450544 520328
rect 450596 520316 450602 520328
rect 477494 520316 477500 520328
rect 450596 520288 477500 520316
rect 450596 520276 450602 520288
rect 477494 520276 477500 520288
rect 477552 520276 477558 520328
rect 353018 520208 353024 520260
rect 353076 520248 353082 520260
rect 357434 520248 357440 520260
rect 353076 520220 357440 520248
rect 353076 520208 353082 520220
rect 357434 520208 357440 520220
rect 357492 520208 357498 520260
rect 401594 520140 401600 520192
rect 401652 520180 401658 520192
rect 403802 520180 403808 520192
rect 401652 520152 403808 520180
rect 401652 520140 401658 520152
rect 403802 520140 403808 520152
rect 403860 520140 403866 520192
rect 322842 519528 322848 519580
rect 322900 519568 322906 519580
rect 324222 519568 324228 519580
rect 322900 519540 324228 519568
rect 322900 519528 322906 519540
rect 324222 519528 324228 519540
rect 324280 519568 324286 519580
rect 355410 519568 355416 519580
rect 324280 519540 355416 519568
rect 324280 519528 324286 519540
rect 355410 519528 355416 519540
rect 355468 519528 355474 519580
rect 321554 519256 321560 519308
rect 321612 519296 321618 519308
rect 323670 519296 323676 519308
rect 321612 519268 323676 519296
rect 321612 519256 321618 519268
rect 323670 519256 323676 519268
rect 323728 519256 323734 519308
rect 454678 518916 454684 518968
rect 454736 518956 454742 518968
rect 478506 518956 478512 518968
rect 454736 518928 478512 518956
rect 454736 518916 454742 518928
rect 478506 518916 478512 518928
rect 478564 518916 478570 518968
rect 513282 518916 513288 518968
rect 513340 518956 513346 518968
rect 531958 518956 531964 518968
rect 513340 518928 531964 518956
rect 513340 518916 513346 518928
rect 531958 518916 531964 518928
rect 532016 518916 532022 518968
rect 321830 518848 321836 518900
rect 321888 518888 321894 518900
rect 325694 518888 325700 518900
rect 321888 518860 325700 518888
rect 321888 518848 321894 518860
rect 325694 518848 325700 518860
rect 325752 518848 325758 518900
rect 345658 518848 345664 518900
rect 345716 518888 345722 518900
rect 357434 518888 357440 518900
rect 345716 518860 357440 518888
rect 345716 518848 345722 518860
rect 357434 518848 357440 518860
rect 357492 518848 357498 518900
rect 322474 517556 322480 517608
rect 322532 517596 322538 517608
rect 350534 517596 350540 517608
rect 322532 517568 350540 517596
rect 322532 517556 322538 517568
rect 350534 517556 350540 517568
rect 350592 517596 350598 517608
rect 356882 517596 356888 517608
rect 350592 517568 356888 517596
rect 350592 517556 350598 517568
rect 356882 517556 356888 517568
rect 356940 517556 356946 517608
rect 466454 517556 466460 517608
rect 466512 517596 466518 517608
rect 477586 517596 477592 517608
rect 466512 517568 477592 517596
rect 466512 517556 466518 517568
rect 477586 517556 477592 517568
rect 477644 517556 477650 517608
rect 254486 517488 254492 517540
rect 254544 517528 254550 517540
rect 274082 517528 274088 517540
rect 254544 517500 274088 517528
rect 254544 517488 254550 517500
rect 274082 517488 274088 517500
rect 274140 517488 274146 517540
rect 326338 517488 326344 517540
rect 326396 517528 326402 517540
rect 357526 517528 357532 517540
rect 326396 517500 357532 517528
rect 326396 517488 326402 517500
rect 357526 517488 357532 517500
rect 357584 517488 357590 517540
rect 436738 517488 436744 517540
rect 436796 517528 436802 517540
rect 477494 517528 477500 517540
rect 436796 517500 477500 517528
rect 436796 517488 436802 517500
rect 477494 517488 477500 517500
rect 477552 517488 477558 517540
rect 321554 517420 321560 517472
rect 321612 517460 321618 517472
rect 323762 517460 323768 517472
rect 321612 517432 323768 517460
rect 321612 517420 321618 517432
rect 323762 517420 323768 517432
rect 323820 517420 323826 517472
rect 341518 517420 341524 517472
rect 341576 517460 341582 517472
rect 357434 517460 357440 517472
rect 341576 517432 357440 517460
rect 341576 517420 341582 517432
rect 357434 517420 357440 517432
rect 357492 517420 357498 517472
rect 477126 517420 477132 517472
rect 477184 517460 477190 517472
rect 478506 517460 478512 517472
rect 477184 517432 478512 517460
rect 477184 517420 477190 517432
rect 478506 517420 478512 517432
rect 478564 517420 478570 517472
rect 322382 516740 322388 516792
rect 322440 516780 322446 516792
rect 322440 516752 335354 516780
rect 322440 516740 322446 516752
rect 335326 516712 335354 516752
rect 356882 516712 356888 516724
rect 335326 516684 356888 516712
rect 356882 516672 356888 516684
rect 356940 516672 356946 516724
rect 322382 516332 322388 516384
rect 322440 516372 322446 516384
rect 322934 516372 322940 516384
rect 322440 516344 322940 516372
rect 322440 516332 322446 516344
rect 322934 516332 322940 516344
rect 322992 516372 322998 516384
rect 325050 516372 325056 516384
rect 322992 516344 325056 516372
rect 322992 516332 322998 516344
rect 325050 516332 325056 516344
rect 325108 516332 325114 516384
rect 513190 516196 513196 516248
rect 513248 516236 513254 516248
rect 526438 516236 526444 516248
rect 513248 516208 526444 516236
rect 513248 516196 513254 516208
rect 526438 516196 526444 516208
rect 526496 516196 526502 516248
rect 402606 516128 402612 516180
rect 402664 516168 402670 516180
rect 405918 516168 405924 516180
rect 402664 516140 405924 516168
rect 402664 516128 402670 516140
rect 405918 516128 405924 516140
rect 405976 516128 405982 516180
rect 513282 516128 513288 516180
rect 513340 516168 513346 516180
rect 536098 516168 536104 516180
rect 513340 516140 536104 516168
rect 513340 516128 513346 516140
rect 536098 516128 536104 516140
rect 536156 516128 536162 516180
rect 321830 516060 321836 516112
rect 321888 516100 321894 516112
rect 342254 516100 342260 516112
rect 321888 516072 342260 516100
rect 321888 516060 321894 516072
rect 342254 516060 342260 516072
rect 342312 516060 342318 516112
rect 401594 516060 401600 516112
rect 401652 516100 401658 516112
rect 403434 516100 403440 516112
rect 401652 516072 403440 516100
rect 401652 516060 401658 516072
rect 403434 516060 403440 516072
rect 403492 516060 403498 516112
rect 513190 516060 513196 516112
rect 513248 516100 513254 516112
rect 520918 516100 520924 516112
rect 513248 516072 520924 516100
rect 513248 516060 513254 516072
rect 520918 516060 520924 516072
rect 520976 516060 520982 516112
rect 322842 515380 322848 515432
rect 322900 515420 322906 515432
rect 324222 515420 324228 515432
rect 322900 515392 324228 515420
rect 322900 515380 322906 515392
rect 324222 515380 324228 515392
rect 324280 515420 324286 515432
rect 329282 515420 329288 515432
rect 324280 515392 329288 515420
rect 324280 515380 324286 515392
rect 329282 515380 329288 515392
rect 329340 515380 329346 515432
rect 342254 515380 342260 515432
rect 342312 515420 342318 515432
rect 343542 515420 343548 515432
rect 342312 515392 343548 515420
rect 342312 515380 342318 515392
rect 343542 515380 343548 515392
rect 343600 515420 343606 515432
rect 353018 515420 353024 515432
rect 343600 515392 353024 515420
rect 343600 515380 343606 515392
rect 353018 515380 353024 515392
rect 353076 515380 353082 515432
rect 358078 514836 358084 514888
rect 358136 514876 358142 514888
rect 359550 514876 359556 514888
rect 358136 514848 359556 514876
rect 358136 514836 358142 514848
rect 359550 514836 359556 514848
rect 359608 514836 359614 514888
rect 331950 514700 331956 514752
rect 332008 514740 332014 514752
rect 357434 514740 357440 514752
rect 332008 514712 357440 514740
rect 332008 514700 332014 514712
rect 357434 514700 357440 514712
rect 357492 514700 357498 514752
rect 322106 514020 322112 514072
rect 322164 514060 322170 514072
rect 332042 514060 332048 514072
rect 322164 514032 332048 514060
rect 322164 514020 322170 514032
rect 332042 514020 332048 514032
rect 332100 514020 332106 514072
rect 460198 513408 460204 513460
rect 460256 513448 460262 513460
rect 477586 513448 477592 513460
rect 460256 513420 477592 513448
rect 460256 513408 460262 513420
rect 477586 513408 477592 513420
rect 477644 513408 477650 513460
rect 322474 513340 322480 513392
rect 322532 513380 322538 513392
rect 355318 513380 355324 513392
rect 322532 513352 355324 513380
rect 322532 513340 322538 513352
rect 355318 513340 355324 513352
rect 355376 513340 355382 513392
rect 441614 513340 441620 513392
rect 441672 513380 441678 513392
rect 477494 513380 477500 513392
rect 441672 513352 477500 513380
rect 441672 513340 441678 513352
rect 477494 513340 477500 513352
rect 477552 513340 477558 513392
rect 320358 513272 320364 513324
rect 320416 513312 320422 513324
rect 355686 513312 355692 513324
rect 320416 513284 355692 513312
rect 320416 513272 320422 513284
rect 355686 513272 355692 513284
rect 355744 513272 355750 513324
rect 358262 513272 358268 513324
rect 358320 513312 358326 513324
rect 359458 513312 359464 513324
rect 358320 513284 359464 513312
rect 358320 513272 358326 513284
rect 359458 513272 359464 513284
rect 359516 513272 359522 513324
rect 412634 513272 412640 513324
rect 412692 513312 412698 513324
rect 477586 513312 477592 513324
rect 412692 513284 477592 513312
rect 412692 513272 412698 513284
rect 477586 513272 477592 513284
rect 477644 513272 477650 513324
rect 329190 513204 329196 513256
rect 329248 513244 329254 513256
rect 357434 513244 357440 513256
rect 329248 513216 357440 513244
rect 329248 513204 329254 513216
rect 357434 513204 357440 513216
rect 357492 513204 357498 513256
rect 402514 513204 402520 513256
rect 402572 513244 402578 513256
rect 405734 513244 405740 513256
rect 402572 513216 405740 513244
rect 402572 513204 402578 513216
rect 405734 513204 405740 513216
rect 405792 513204 405798 513256
rect 322106 512592 322112 512644
rect 322164 512632 322170 512644
rect 357158 512632 357164 512644
rect 322164 512604 357164 512632
rect 322164 512592 322170 512604
rect 357158 512592 357164 512604
rect 357216 512592 357222 512644
rect 340230 511912 340236 511964
rect 340288 511952 340294 511964
rect 357434 511952 357440 511964
rect 340288 511924 357440 511952
rect 340288 511912 340294 511924
rect 357434 511912 357440 511924
rect 357492 511912 357498 511964
rect 321554 511232 321560 511284
rect 321612 511272 321618 511284
rect 336642 511272 336648 511284
rect 321612 511244 336648 511272
rect 321612 511232 321618 511244
rect 336642 511232 336648 511244
rect 336700 511272 336706 511284
rect 356974 511272 356980 511284
rect 336700 511244 356980 511272
rect 336700 511232 336706 511244
rect 356974 511232 356980 511244
rect 357032 511232 357038 511284
rect 320358 510824 320364 510876
rect 320416 510864 320422 510876
rect 320634 510864 320640 510876
rect 320416 510836 320640 510864
rect 320416 510824 320422 510836
rect 320634 510824 320640 510836
rect 320692 510864 320698 510876
rect 327902 510864 327908 510876
rect 320692 510836 327908 510864
rect 320692 510824 320698 510836
rect 327902 510824 327908 510836
rect 327960 510824 327966 510876
rect 254394 510620 254400 510672
rect 254452 510660 254458 510672
rect 271322 510660 271328 510672
rect 254452 510632 271328 510660
rect 254452 510620 254458 510632
rect 271322 510620 271328 510632
rect 271380 510620 271386 510672
rect 402882 510620 402888 510672
rect 402940 510660 402946 510672
rect 451274 510660 451280 510672
rect 402940 510632 451280 510660
rect 402940 510620 402946 510632
rect 451274 510620 451280 510632
rect 451332 510620 451338 510672
rect 462958 510620 462964 510672
rect 463016 510660 463022 510672
rect 477586 510660 477592 510672
rect 463016 510632 477592 510660
rect 463016 510620 463022 510632
rect 477586 510620 477592 510632
rect 477644 510620 477650 510672
rect 513282 510620 513288 510672
rect 513340 510660 513346 510672
rect 544378 510660 544384 510672
rect 513340 510632 544384 510660
rect 513340 510620 513346 510632
rect 544378 510620 544384 510632
rect 544436 510620 544442 510672
rect 320082 510552 320088 510604
rect 320140 510592 320146 510604
rect 355594 510592 355600 510604
rect 320140 510564 355600 510592
rect 320140 510552 320146 510564
rect 355594 510552 355600 510564
rect 355652 510552 355658 510604
rect 462314 510552 462320 510604
rect 462372 510592 462378 510604
rect 477494 510592 477500 510604
rect 462372 510564 477500 510592
rect 462372 510552 462378 510564
rect 477494 510552 477500 510564
rect 477552 510552 477558 510604
rect 320450 510484 320456 510536
rect 320508 510524 320514 510536
rect 333330 510524 333336 510536
rect 320508 510496 333336 510524
rect 320508 510484 320514 510496
rect 333330 510484 333336 510496
rect 333388 510484 333394 510536
rect 337562 510484 337568 510536
rect 337620 510524 337626 510536
rect 357434 510524 357440 510536
rect 337620 510496 357440 510524
rect 337620 510484 337626 510496
rect 357434 510484 357440 510496
rect 357492 510484 357498 510536
rect 324222 509872 324228 509924
rect 324280 509912 324286 509924
rect 350074 509912 350080 509924
rect 324280 509884 350080 509912
rect 324280 509872 324286 509884
rect 350074 509872 350080 509884
rect 350132 509872 350138 509924
rect 402882 509328 402888 509380
rect 402940 509368 402946 509380
rect 404906 509368 404912 509380
rect 402940 509340 404912 509368
rect 402940 509328 402946 509340
rect 404906 509328 404912 509340
rect 404964 509368 404970 509380
rect 445018 509368 445024 509380
rect 404964 509340 445024 509368
rect 404964 509328 404970 509340
rect 445018 509328 445024 509340
rect 445076 509328 445082 509380
rect 422938 509260 422944 509312
rect 422996 509300 423002 509312
rect 477494 509300 477500 509312
rect 422996 509272 477500 509300
rect 422996 509260 423002 509272
rect 477494 509260 477500 509272
rect 477552 509260 477558 509312
rect 513282 509260 513288 509312
rect 513340 509300 513346 509312
rect 522298 509300 522304 509312
rect 513340 509272 522304 509300
rect 513340 509260 513346 509272
rect 522298 509260 522304 509272
rect 522356 509260 522362 509312
rect 320174 509192 320180 509244
rect 320232 509232 320238 509244
rect 353202 509232 353208 509244
rect 320232 509204 353208 509232
rect 320232 509192 320238 509204
rect 353202 509192 353208 509204
rect 353260 509192 353266 509244
rect 342898 509124 342904 509176
rect 342956 509164 342962 509176
rect 357526 509164 357532 509176
rect 342956 509136 357532 509164
rect 342956 509124 342962 509136
rect 357526 509124 357532 509136
rect 357584 509124 357590 509176
rect 347038 509056 347044 509108
rect 347096 509096 347102 509108
rect 357434 509096 357440 509108
rect 347096 509068 357440 509096
rect 347096 509056 347102 509068
rect 357434 509056 357440 509068
rect 357492 509056 357498 509108
rect 478782 508444 478788 508496
rect 478840 508484 478846 508496
rect 479518 508484 479524 508496
rect 478840 508456 479524 508484
rect 478840 508444 478846 508456
rect 479518 508444 479524 508456
rect 479576 508444 479582 508496
rect 319070 508240 319076 508292
rect 319128 508280 319134 508292
rect 319346 508280 319352 508292
rect 319128 508252 319352 508280
rect 319128 508240 319134 508252
rect 319346 508240 319352 508252
rect 319404 508240 319410 508292
rect 50798 507832 50804 507884
rect 50856 507872 50862 507884
rect 51166 507872 51172 507884
rect 50856 507844 51172 507872
rect 50856 507832 50862 507844
rect 51166 507832 51172 507844
rect 51224 507832 51230 507884
rect 319070 507832 319076 507884
rect 319128 507872 319134 507884
rect 357158 507872 357164 507884
rect 319128 507844 357164 507872
rect 319128 507832 319134 507844
rect 357158 507832 357164 507844
rect 357216 507832 357222 507884
rect 358722 507832 358728 507884
rect 358780 507872 358786 507884
rect 359734 507872 359740 507884
rect 358780 507844 359740 507872
rect 358780 507832 358786 507844
rect 359734 507832 359740 507844
rect 359792 507832 359798 507884
rect 320358 507764 320364 507816
rect 320416 507804 320422 507816
rect 355502 507804 355508 507816
rect 320416 507776 355508 507804
rect 320416 507764 320422 507776
rect 355502 507764 355508 507776
rect 355560 507764 355566 507816
rect 334618 507696 334624 507748
rect 334676 507736 334682 507748
rect 357434 507736 357440 507748
rect 334676 507708 357440 507736
rect 334676 507696 334682 507708
rect 357434 507696 357440 507708
rect 357492 507696 357498 507748
rect 320082 507628 320088 507680
rect 320140 507668 320146 507680
rect 345842 507668 345848 507680
rect 320140 507640 345848 507668
rect 320140 507628 320146 507640
rect 345842 507628 345848 507640
rect 345900 507628 345906 507680
rect 318978 506472 318984 506524
rect 319036 506512 319042 506524
rect 320082 506512 320088 506524
rect 319036 506484 320088 506512
rect 319036 506472 319042 506484
rect 320082 506472 320088 506484
rect 320140 506472 320146 506524
rect 320174 506404 320180 506456
rect 320232 506444 320238 506456
rect 345750 506444 345756 506456
rect 320232 506416 345756 506444
rect 320232 506404 320238 506416
rect 345750 506404 345756 506416
rect 345808 506404 345814 506456
rect 347130 506404 347136 506456
rect 347188 506444 347194 506456
rect 357434 506444 357440 506456
rect 347188 506416 357440 506444
rect 347188 506404 347194 506416
rect 357434 506404 357440 506416
rect 357492 506404 357498 506456
rect 402238 506404 402244 506456
rect 402296 506444 402302 506456
rect 404814 506444 404820 506456
rect 402296 506416 404820 506444
rect 402296 506404 402302 506416
rect 404814 506404 404820 506416
rect 404872 506404 404878 506456
rect 349982 506336 349988 506388
rect 350040 506376 350046 506388
rect 357526 506376 357532 506388
rect 350040 506348 357532 506376
rect 350040 506336 350046 506348
rect 357526 506336 357532 506348
rect 357584 506336 357590 506388
rect 319346 505724 319352 505776
rect 319404 505764 319410 505776
rect 325510 505764 325516 505776
rect 319404 505736 325516 505764
rect 319404 505724 319410 505736
rect 325510 505724 325516 505736
rect 325568 505764 325574 505776
rect 356606 505764 356612 505776
rect 325568 505736 356612 505764
rect 325568 505724 325574 505736
rect 356606 505724 356612 505736
rect 356664 505724 356670 505776
rect 318886 505520 318892 505572
rect 318944 505560 318950 505572
rect 319346 505560 319352 505572
rect 318944 505532 319352 505560
rect 318944 505520 318950 505532
rect 319346 505520 319352 505532
rect 319404 505520 319410 505572
rect 472710 505520 472716 505572
rect 472768 505560 472774 505572
rect 477494 505560 477500 505572
rect 472768 505532 477500 505560
rect 472768 505520 472774 505532
rect 477494 505520 477500 505532
rect 477552 505520 477558 505572
rect 254302 505112 254308 505164
rect 254360 505152 254366 505164
rect 275462 505152 275468 505164
rect 254360 505124 275468 505152
rect 254360 505112 254366 505124
rect 275462 505112 275468 505124
rect 275520 505112 275526 505164
rect 320174 505112 320180 505164
rect 320232 505152 320238 505164
rect 320726 505152 320732 505164
rect 320232 505124 320732 505152
rect 320232 505112 320238 505124
rect 320726 505112 320732 505124
rect 320784 505112 320790 505164
rect 340874 505112 340880 505164
rect 340932 505152 340938 505164
rect 342162 505152 342168 505164
rect 340932 505124 342168 505152
rect 340932 505112 340938 505124
rect 342162 505112 342168 505124
rect 342220 505152 342226 505164
rect 359734 505152 359740 505164
rect 342220 505124 359740 505152
rect 342220 505112 342226 505124
rect 359734 505112 359740 505124
rect 359792 505112 359798 505164
rect 404998 505112 405004 505164
rect 405056 505152 405062 505164
rect 477494 505152 477500 505164
rect 405056 505124 477500 505152
rect 405056 505112 405062 505124
rect 477494 505112 477500 505124
rect 477552 505112 477558 505164
rect 327718 505044 327724 505096
rect 327776 505084 327782 505096
rect 357434 505084 357440 505096
rect 327776 505056 357440 505084
rect 327776 505044 327782 505056
rect 357434 505044 357440 505056
rect 357492 505044 357498 505096
rect 320082 504976 320088 505028
rect 320140 505016 320146 505028
rect 340874 505016 340880 505028
rect 320140 504988 340880 505016
rect 320140 504976 320146 504988
rect 340874 504976 340880 504988
rect 340932 504976 340938 505028
rect 322382 504160 322388 504212
rect 322440 504200 322446 504212
rect 326338 504200 326344 504212
rect 322440 504172 326344 504200
rect 322440 504160 322446 504172
rect 326338 504160 326344 504172
rect 326396 504160 326402 504212
rect 436830 503752 436836 503804
rect 436888 503792 436894 503804
rect 477586 503792 477592 503804
rect 436888 503764 477592 503792
rect 436888 503752 436894 503764
rect 477586 503752 477592 503764
rect 477644 503752 477650 503804
rect 400858 503684 400864 503736
rect 400916 503724 400922 503736
rect 477494 503724 477500 503736
rect 400916 503696 477500 503724
rect 400916 503684 400922 503696
rect 477494 503684 477500 503696
rect 477552 503684 477558 503736
rect 513282 503684 513288 503736
rect 513340 503724 513346 503736
rect 530578 503724 530584 503736
rect 513340 503696 530584 503724
rect 513340 503684 513346 503696
rect 530578 503684 530584 503696
rect 530636 503684 530642 503736
rect 320174 503616 320180 503668
rect 320232 503656 320238 503668
rect 325602 503656 325608 503668
rect 320232 503628 325608 503656
rect 320232 503616 320238 503628
rect 325602 503616 325608 503628
rect 325660 503656 325666 503668
rect 357434 503656 357440 503668
rect 325660 503628 357440 503656
rect 325660 503616 325666 503628
rect 357434 503616 357440 503628
rect 357492 503616 357498 503668
rect 401686 503616 401692 503668
rect 401744 503656 401750 503668
rect 405826 503656 405832 503668
rect 401744 503628 405832 503656
rect 401744 503616 401750 503628
rect 405826 503616 405832 503628
rect 405884 503616 405890 503668
rect 322382 503548 322388 503600
rect 322440 503588 322446 503600
rect 348418 503588 348424 503600
rect 322440 503560 348424 503588
rect 322440 503548 322446 503560
rect 348418 503548 348424 503560
rect 348476 503548 348482 503600
rect 478506 502596 478512 502648
rect 478564 502636 478570 502648
rect 478782 502636 478788 502648
rect 478564 502608 478788 502636
rect 478564 502596 478570 502608
rect 478782 502596 478788 502608
rect 478840 502596 478846 502648
rect 322382 502324 322388 502376
rect 322440 502364 322446 502376
rect 355502 502364 355508 502376
rect 322440 502336 355508 502364
rect 322440 502324 322446 502336
rect 355502 502324 355508 502336
rect 355560 502324 355566 502376
rect 440878 502324 440884 502376
rect 440936 502364 440942 502376
rect 477494 502364 477500 502376
rect 440936 502336 477500 502364
rect 440936 502324 440942 502336
rect 477494 502324 477500 502336
rect 477552 502324 477558 502376
rect 513282 502324 513288 502376
rect 513340 502364 513346 502376
rect 545758 502364 545764 502376
rect 513340 502336 545764 502364
rect 513340 502324 513346 502336
rect 545758 502324 545764 502336
rect 545816 502324 545822 502376
rect 337378 502256 337384 502308
rect 337436 502296 337442 502308
rect 357434 502296 357440 502308
rect 337436 502268 357440 502296
rect 337436 502256 337442 502268
rect 357434 502256 357440 502268
rect 357492 502256 357498 502308
rect 402238 500964 402244 501016
rect 402296 501004 402302 501016
rect 477494 501004 477500 501016
rect 402296 500976 477500 501004
rect 402296 500964 402302 500976
rect 477494 500964 477500 500976
rect 477552 500964 477558 501016
rect 352558 500896 352564 500948
rect 352616 500936 352622 500948
rect 399478 500936 399484 500948
rect 352616 500908 399484 500936
rect 352616 500896 352622 500908
rect 399478 500896 399484 500908
rect 399536 500896 399542 500948
rect 478598 500896 478604 500948
rect 478656 500936 478662 500948
rect 510706 500936 510712 500948
rect 478656 500908 510712 500936
rect 478656 500896 478662 500908
rect 510706 500896 510712 500908
rect 510764 500896 510770 500948
rect 353110 500828 353116 500880
rect 353168 500868 353174 500880
rect 402054 500868 402060 500880
rect 353168 500840 402060 500868
rect 353168 500828 353174 500840
rect 402054 500828 402060 500840
rect 402112 500828 402118 500880
rect 358354 500760 358360 500812
rect 358412 500800 358418 500812
rect 359366 500800 359372 500812
rect 358412 500772 359372 500800
rect 358412 500760 358418 500772
rect 359366 500760 359372 500772
rect 359424 500760 359430 500812
rect 510706 500760 510712 500812
rect 510764 500800 510770 500812
rect 510982 500800 510988 500812
rect 510764 500772 510988 500800
rect 510764 500760 510770 500772
rect 510982 500760 510988 500772
rect 511040 500760 511046 500812
rect 510982 500624 510988 500676
rect 511040 500664 511046 500676
rect 511258 500664 511264 500676
rect 511040 500636 511264 500664
rect 511040 500624 511046 500636
rect 511258 500624 511264 500636
rect 511316 500624 511322 500676
rect 296622 500352 296628 500404
rect 296680 500392 296686 500404
rect 321738 500392 321744 500404
rect 296680 500364 321744 500392
rect 296680 500352 296686 500364
rect 321738 500352 321744 500364
rect 321796 500352 321802 500404
rect 295242 500284 295248 500336
rect 295300 500324 295306 500336
rect 321646 500324 321652 500336
rect 295300 500296 321652 500324
rect 295300 500284 295306 500296
rect 321646 500284 321652 500296
rect 321704 500284 321710 500336
rect 292758 500216 292764 500268
rect 292816 500256 292822 500268
rect 320634 500256 320640 500268
rect 292816 500228 320640 500256
rect 292816 500216 292822 500228
rect 320634 500216 320640 500228
rect 320692 500216 320698 500268
rect 322198 500216 322204 500268
rect 322256 500256 322262 500268
rect 322256 500228 354674 500256
rect 322256 500216 322262 500228
rect 354646 499984 354674 500228
rect 360838 499984 360844 499996
rect 354646 499956 360844 499984
rect 360838 499944 360844 499956
rect 360896 499944 360902 499996
rect 254210 499876 254216 499928
rect 254268 499916 254274 499928
rect 257430 499916 257436 499928
rect 254268 499888 257436 499916
rect 254268 499876 254274 499888
rect 257430 499876 257436 499888
rect 257488 499876 257494 499928
rect 401870 499536 401876 499588
rect 401928 499576 401934 499588
rect 433334 499576 433340 499588
rect 401928 499548 433340 499576
rect 401928 499536 401934 499548
rect 433334 499536 433340 499548
rect 433392 499536 433398 499588
rect 468570 499536 468576 499588
rect 468628 499576 468634 499588
rect 477494 499576 477500 499588
rect 468628 499548 477500 499576
rect 468628 499536 468634 499548
rect 477494 499536 477500 499548
rect 477552 499536 477558 499588
rect 355962 499468 355968 499520
rect 356020 499508 356026 499520
rect 364518 499508 364524 499520
rect 356020 499480 364524 499508
rect 356020 499468 356026 499480
rect 364518 499468 364524 499480
rect 364576 499468 364582 499520
rect 394142 499468 394148 499520
rect 394200 499508 394206 499520
rect 403710 499508 403716 499520
rect 394200 499480 403716 499508
rect 394200 499468 394206 499480
rect 403710 499468 403716 499480
rect 403768 499468 403774 499520
rect 478782 499468 478788 499520
rect 478840 499508 478846 499520
rect 482370 499508 482376 499520
rect 478840 499480 482376 499508
rect 478840 499468 478846 499480
rect 482370 499468 482376 499480
rect 482428 499468 482434 499520
rect 373534 499400 373540 499452
rect 373592 499440 373598 499452
rect 471238 499440 471244 499452
rect 373592 499412 471244 499440
rect 373592 499400 373598 499412
rect 471238 499400 471244 499412
rect 471296 499400 471302 499452
rect 487798 499400 487804 499452
rect 487856 499440 487862 499452
rect 525150 499440 525156 499452
rect 487856 499412 525156 499440
rect 487856 499400 487862 499412
rect 525150 499400 525156 499412
rect 525208 499400 525214 499452
rect 322290 499332 322296 499384
rect 322348 499372 322354 499384
rect 400766 499372 400772 499384
rect 322348 499344 400772 499372
rect 322348 499332 322354 499344
rect 400766 499332 400772 499344
rect 400824 499332 400830 499384
rect 477034 499332 477040 499384
rect 477092 499372 477098 499384
rect 499298 499372 499304 499384
rect 477092 499344 499304 499372
rect 477092 499332 477098 499344
rect 499298 499332 499304 499344
rect 499356 499332 499362 499384
rect 353018 499264 353024 499316
rect 353076 499304 353082 499316
rect 398006 499304 398012 499316
rect 353076 499276 398012 499304
rect 353076 499264 353082 499276
rect 398006 499264 398012 499276
rect 398064 499264 398070 499316
rect 492306 499264 492312 499316
rect 492364 499304 492370 499316
rect 511350 499304 511356 499316
rect 492364 499276 511356 499304
rect 492364 499264 492370 499276
rect 511350 499264 511356 499276
rect 511408 499264 511414 499316
rect 359826 499196 359832 499248
rect 359884 499236 359890 499248
rect 401686 499236 401692 499248
rect 359884 499208 401692 499236
rect 359884 499196 359890 499208
rect 401686 499196 401692 499208
rect 401744 499196 401750 499248
rect 359734 499128 359740 499180
rect 359792 499168 359798 499180
rect 401594 499168 401600 499180
rect 359792 499140 401600 499168
rect 359792 499128 359798 499140
rect 401594 499128 401600 499140
rect 401652 499128 401658 499180
rect 359918 499060 359924 499112
rect 359976 499100 359982 499112
rect 401962 499100 401968 499112
rect 359976 499072 401968 499100
rect 359976 499060 359982 499072
rect 401962 499060 401968 499072
rect 402020 499060 402026 499112
rect 357066 498992 357072 499044
rect 357124 499032 357130 499044
rect 397362 499032 397368 499044
rect 357124 499004 397368 499032
rect 357124 498992 357130 499004
rect 397362 498992 397368 499004
rect 397420 498992 397426 499044
rect 356606 498924 356612 498976
rect 356664 498964 356670 498976
rect 381906 498964 381912 498976
rect 356664 498936 381912 498964
rect 356664 498924 356670 498936
rect 381906 498924 381912 498936
rect 381964 498924 381970 498976
rect 323670 498856 323676 498908
rect 323728 498896 323734 498908
rect 353386 498896 353392 498908
rect 323728 498868 353392 498896
rect 323728 498856 323734 498868
rect 353386 498856 353392 498868
rect 353444 498896 353450 498908
rect 367738 498896 367744 498908
rect 353444 498868 367744 498896
rect 353444 498856 353450 498868
rect 367738 498856 367744 498868
rect 367796 498856 367802 498908
rect 254578 498788 254584 498840
rect 254636 498828 254642 498840
rect 282178 498828 282184 498840
rect 254636 498800 282184 498828
rect 254636 498788 254642 498800
rect 282178 498788 282184 498800
rect 282236 498788 282242 498840
rect 322474 498788 322480 498840
rect 322532 498828 322538 498840
rect 362954 498828 362960 498840
rect 322532 498800 362960 498828
rect 322532 498788 322538 498800
rect 362954 498788 362960 498800
rect 363012 498788 363018 498840
rect 508498 498788 508504 498840
rect 508556 498828 508562 498840
rect 511994 498828 512000 498840
rect 508556 498800 512000 498828
rect 508556 498788 508562 498800
rect 511994 498788 512000 498800
rect 512052 498788 512058 498840
rect 356974 498720 356980 498772
rect 357032 498760 357038 498772
rect 389634 498760 389640 498772
rect 357032 498732 389640 498760
rect 357032 498720 357038 498732
rect 389634 498720 389640 498732
rect 389692 498720 389698 498772
rect 479242 498720 479248 498772
rect 479300 498760 479306 498772
rect 481634 498760 481640 498772
rect 479300 498732 481640 498760
rect 479300 498720 479306 498732
rect 481634 498720 481640 498732
rect 481692 498720 481698 498772
rect 375466 498652 375472 498704
rect 375524 498692 375530 498704
rect 580350 498692 580356 498704
rect 375524 498664 580356 498692
rect 375524 498652 375530 498664
rect 580350 498652 580356 498664
rect 580408 498652 580414 498704
rect 324958 498584 324964 498636
rect 325016 498624 325022 498636
rect 378042 498624 378048 498636
rect 325016 498596 378048 498624
rect 325016 498584 325022 498596
rect 378042 498584 378048 498596
rect 378100 498584 378106 498636
rect 352558 498176 352564 498228
rect 352616 498216 352622 498228
rect 353018 498216 353024 498228
rect 352616 498188 353024 498216
rect 352616 498176 352622 498188
rect 353018 498176 353024 498188
rect 353076 498176 353082 498228
rect 478414 498176 478420 498228
rect 478472 498216 478478 498228
rect 480898 498216 480904 498228
rect 478472 498188 480904 498216
rect 478472 498176 478478 498188
rect 480898 498176 480904 498188
rect 480956 498176 480962 498228
rect 352834 498108 352840 498160
rect 352892 498148 352898 498160
rect 355318 498148 355324 498160
rect 352892 498120 355324 498148
rect 352892 498108 352898 498120
rect 355318 498108 355324 498120
rect 355376 498108 355382 498160
rect 355410 498108 355416 498160
rect 355468 498148 355474 498160
rect 361298 498148 361304 498160
rect 355468 498120 361304 498148
rect 355468 498108 355474 498120
rect 361298 498108 361304 498120
rect 361356 498108 361362 498160
rect 399294 498108 399300 498160
rect 399352 498148 399358 498160
rect 403894 498148 403900 498160
rect 399352 498120 403900 498148
rect 399352 498108 399358 498120
rect 403894 498108 403900 498120
rect 403952 498108 403958 498160
rect 475654 498108 475660 498160
rect 475712 498148 475718 498160
rect 484486 498148 484492 498160
rect 475712 498120 484492 498148
rect 475712 498108 475718 498120
rect 484486 498108 484492 498120
rect 484544 498108 484550 498160
rect 491018 498108 491024 498160
rect 491076 498148 491082 498160
rect 521654 498148 521660 498160
rect 491076 498120 521660 498148
rect 491076 498108 491082 498120
rect 521654 498108 521660 498120
rect 521712 498108 521718 498160
rect 357342 498040 357348 498092
rect 357400 498080 357406 498092
rect 370958 498080 370964 498092
rect 357400 498052 370964 498080
rect 357400 498040 357406 498052
rect 370958 498040 370964 498052
rect 371016 498040 371022 498092
rect 396718 498040 396724 498092
rect 396776 498080 396782 498092
rect 405182 498080 405188 498092
rect 396776 498052 405188 498080
rect 396776 498040 396782 498052
rect 405182 498040 405188 498052
rect 405240 498040 405246 498092
rect 473998 498040 474004 498092
rect 474056 498080 474062 498092
rect 503162 498080 503168 498092
rect 474056 498052 503168 498080
rect 474056 498040 474062 498052
rect 503162 498040 503168 498052
rect 503220 498040 503226 498092
rect 357250 497972 357256 498024
rect 357308 498012 357314 498024
rect 367094 498012 367100 498024
rect 357308 497984 367100 498012
rect 357308 497972 357314 497984
rect 367094 497972 367100 497984
rect 367152 497972 367158 498024
rect 388346 497972 388352 498024
rect 388404 498012 388410 498024
rect 405274 498012 405280 498024
rect 388404 497984 405280 498012
rect 388404 497972 388410 497984
rect 405274 497972 405280 497984
rect 405332 497972 405338 498024
rect 475838 497972 475844 498024
rect 475896 498012 475902 498024
rect 502518 498012 502524 498024
rect 475896 497984 502524 498012
rect 475896 497972 475902 497984
rect 502518 497972 502524 497984
rect 502576 497972 502582 498024
rect 294598 497904 294604 497956
rect 294656 497944 294662 497956
rect 316034 497944 316040 497956
rect 294656 497916 316040 497944
rect 294656 497904 294662 497916
rect 316034 497904 316040 497916
rect 316092 497904 316098 497956
rect 349798 497904 349804 497956
rect 349856 497944 349862 497956
rect 379330 497944 379336 497956
rect 349856 497916 379336 497944
rect 349856 497904 349862 497916
rect 379330 497904 379336 497916
rect 379388 497904 379394 497956
rect 477218 497904 477224 497956
rect 477276 497944 477282 497956
rect 496722 497944 496728 497956
rect 477276 497916 496728 497944
rect 477276 497904 477282 497916
rect 496722 497904 496728 497916
rect 496780 497904 496786 497956
rect 291930 497836 291936 497888
rect 291988 497876 291994 497888
rect 315114 497876 315120 497888
rect 291988 497848 315120 497876
rect 291988 497836 291994 497848
rect 315114 497836 315120 497848
rect 315172 497836 315178 497888
rect 352742 497836 352748 497888
rect 352800 497876 352806 497888
rect 379974 497876 379980 497888
rect 352800 497848 379980 497876
rect 352800 497836 352806 497848
rect 379974 497836 379980 497848
rect 380032 497836 380038 497888
rect 494790 497836 494796 497888
rect 494848 497876 494854 497888
rect 510246 497876 510252 497888
rect 494848 497848 510252 497876
rect 494848 497836 494854 497848
rect 510246 497836 510252 497848
rect 510304 497836 510310 497888
rect 290458 497768 290464 497820
rect 290516 497808 290522 497820
rect 327718 497808 327724 497820
rect 290516 497780 327724 497808
rect 290516 497768 290522 497780
rect 327718 497768 327724 497780
rect 327776 497768 327782 497820
rect 352926 497768 352932 497820
rect 352984 497808 352990 497820
rect 366450 497808 366456 497820
rect 352984 497780 366456 497808
rect 352984 497768 352990 497780
rect 366450 497768 366456 497780
rect 366508 497768 366514 497820
rect 470594 497768 470600 497820
rect 470652 497808 470658 497820
rect 485130 497808 485136 497820
rect 470652 497780 485136 497808
rect 470652 497768 470658 497780
rect 485130 497768 485136 497780
rect 485188 497768 485194 497820
rect 258718 497700 258724 497752
rect 258776 497740 258782 497752
rect 301866 497740 301872 497752
rect 258776 497712 301872 497740
rect 258776 497700 258782 497712
rect 301866 497700 301872 497712
rect 301924 497700 301930 497752
rect 355318 497700 355324 497752
rect 355376 497740 355382 497752
rect 363230 497740 363236 497752
rect 355376 497712 363236 497740
rect 355376 497700 355382 497712
rect 363230 497700 363236 497712
rect 363288 497700 363294 497752
rect 260282 497632 260288 497684
rect 260340 497672 260346 497684
rect 316586 497672 316592 497684
rect 260340 497644 316592 497672
rect 260340 497632 260346 497644
rect 316586 497632 316592 497644
rect 316644 497632 316650 497684
rect 351362 497632 351368 497684
rect 351420 497672 351426 497684
rect 394786 497672 394792 497684
rect 351420 497644 394792 497672
rect 351420 497632 351426 497644
rect 394786 497632 394792 497644
rect 394844 497632 394850 497684
rect 427814 497632 427820 497684
rect 427872 497672 427878 497684
rect 493502 497672 493508 497684
rect 427872 497644 493508 497672
rect 427872 497632 427878 497644
rect 493502 497632 493508 497644
rect 493560 497632 493566 497684
rect 257614 497564 257620 497616
rect 257672 497604 257678 497616
rect 317414 497604 317420 497616
rect 257672 497576 317420 497604
rect 257672 497564 257678 497576
rect 317414 497564 317420 497576
rect 317472 497564 317478 497616
rect 352650 497564 352656 497616
rect 352708 497604 352714 497616
rect 372246 497604 372252 497616
rect 352708 497576 372252 497604
rect 352708 497564 352714 497576
rect 372246 497564 372252 497576
rect 372304 497564 372310 497616
rect 459554 497564 459560 497616
rect 459612 497604 459618 497616
rect 505738 497604 505744 497616
rect 459612 497576 505744 497604
rect 459612 497564 459618 497576
rect 505738 497564 505744 497576
rect 505796 497564 505802 497616
rect 254670 497496 254676 497548
rect 254728 497536 254734 497548
rect 314654 497536 314660 497548
rect 254728 497508 314660 497536
rect 254728 497496 254734 497508
rect 314654 497496 314660 497508
rect 314712 497496 314718 497548
rect 414014 497496 414020 497548
rect 414072 497536 414078 497548
rect 492858 497536 492864 497548
rect 414072 497508 492864 497536
rect 414072 497496 414078 497508
rect 492858 497496 492864 497508
rect 492916 497496 492922 497548
rect 296530 497428 296536 497480
rect 296588 497468 296594 497480
rect 487062 497468 487068 497480
rect 296588 497440 487068 497468
rect 296588 497428 296594 497440
rect 487062 497428 487068 497440
rect 487120 497428 487126 497480
rect 493410 497428 493416 497480
rect 493468 497468 493474 497480
rect 507026 497468 507032 497480
rect 493468 497440 507032 497468
rect 493468 497428 493474 497440
rect 507026 497428 507032 497440
rect 507084 497428 507090 497480
rect 359366 497360 359372 497412
rect 359424 497400 359430 497412
rect 481910 497400 481916 497412
rect 359424 497372 481916 497400
rect 359424 497360 359430 497372
rect 481910 497360 481916 497372
rect 481968 497360 481974 497412
rect 354122 497292 354128 497344
rect 354180 497332 354186 497344
rect 383838 497332 383844 497344
rect 354180 497304 383844 497332
rect 354180 497292 354186 497304
rect 383838 497292 383844 497304
rect 383896 497292 383902 497344
rect 496170 496952 496176 497004
rect 496228 496992 496234 497004
rect 501874 496992 501880 497004
rect 496228 496964 501880 496992
rect 496228 496952 496234 496964
rect 501874 496952 501880 496964
rect 501932 496952 501938 497004
rect 494698 496884 494704 496936
rect 494756 496924 494762 496936
rect 498010 496924 498016 496936
rect 494756 496896 498016 496924
rect 494756 496884 494762 496896
rect 498010 496884 498016 496896
rect 498068 496884 498074 496936
rect 502334 496884 502340 496936
rect 502392 496924 502398 496936
rect 509694 496924 509700 496936
rect 502392 496896 509700 496924
rect 502392 496884 502398 496896
rect 509694 496884 509700 496896
rect 509752 496884 509758 496936
rect 284570 496816 284576 496868
rect 284628 496856 284634 496868
rect 286318 496856 286324 496868
rect 284628 496828 286324 496856
rect 284628 496816 284634 496828
rect 286318 496816 286324 496828
rect 286376 496816 286382 496868
rect 299842 496816 299848 496868
rect 299900 496856 299906 496868
rect 305546 496856 305552 496868
rect 299900 496828 305552 496856
rect 299900 496816 299906 496828
rect 305546 496816 305552 496828
rect 305604 496816 305610 496868
rect 381538 496816 381544 496868
rect 381596 496856 381602 496868
rect 384482 496856 384488 496868
rect 381596 496828 384488 496856
rect 381596 496816 381602 496828
rect 384482 496816 384488 496828
rect 384540 496816 384546 496868
rect 485038 496816 485044 496868
rect 485096 496856 485102 496868
rect 488350 496856 488356 496868
rect 485096 496828 488356 496856
rect 485096 496816 485102 496828
rect 488350 496816 488356 496828
rect 488408 496816 488414 496868
rect 493318 496816 493324 496868
rect 493376 496856 493382 496868
rect 494146 496856 494152 496868
rect 493376 496828 494152 496856
rect 493376 496816 493382 496828
rect 494146 496816 494152 496828
rect 494204 496816 494210 496868
rect 496078 496816 496084 496868
rect 496136 496856 496142 496868
rect 498654 496856 498660 496868
rect 496136 496828 498660 496856
rect 496136 496816 496142 496828
rect 498654 496816 498660 496828
rect 498712 496816 498718 496868
rect 502978 496816 502984 496868
rect 503036 496856 503042 496868
rect 503806 496856 503812 496868
rect 503036 496828 503812 496856
rect 503036 496816 503042 496828
rect 503806 496816 503812 496828
rect 503864 496816 503870 496868
rect 358170 496748 358176 496800
rect 358228 496788 358234 496800
rect 366358 496788 366364 496800
rect 358228 496760 366364 496788
rect 358228 496748 358234 496760
rect 366358 496748 366364 496760
rect 366416 496748 366422 496800
rect 478230 496748 478236 496800
rect 478288 496788 478294 496800
rect 482278 496788 482284 496800
rect 478288 496760 482284 496788
rect 478288 496748 478294 496760
rect 482278 496748 482284 496760
rect 482336 496748 482342 496800
rect 294138 496680 294144 496732
rect 294196 496720 294202 496732
rect 295978 496720 295984 496732
rect 294196 496692 295984 496720
rect 294196 496680 294202 496692
rect 295978 496680 295984 496692
rect 296036 496680 296042 496732
rect 479150 496204 479156 496256
rect 479208 496244 479214 496256
rect 488626 496244 488632 496256
rect 479208 496216 488632 496244
rect 479208 496204 479214 496216
rect 488626 496204 488632 496216
rect 488684 496204 488690 496256
rect 278774 496136 278780 496188
rect 278832 496176 278838 496188
rect 320542 496176 320548 496188
rect 278832 496148 320548 496176
rect 278832 496136 278838 496148
rect 320542 496136 320548 496148
rect 320600 496136 320606 496188
rect 479702 496176 479708 496188
rect 470566 496148 479708 496176
rect 264974 496068 264980 496120
rect 265032 496108 265038 496120
rect 320726 496108 320732 496120
rect 265032 496080 320732 496108
rect 265032 496068 265038 496080
rect 320726 496068 320732 496080
rect 320784 496068 320790 496120
rect 367094 496068 367100 496120
rect 367152 496108 367158 496120
rect 470566 496108 470594 496148
rect 479702 496136 479708 496148
rect 479760 496136 479766 496188
rect 495526 496136 495532 496188
rect 495584 496176 495590 496188
rect 552658 496176 552664 496188
rect 495584 496148 552664 496176
rect 495584 496136 495590 496148
rect 552658 496136 552664 496148
rect 552716 496136 552722 496188
rect 367152 496080 470594 496108
rect 367152 496068 367158 496080
rect 479334 496068 479340 496120
rect 479392 496108 479398 496120
rect 547874 496108 547880 496120
rect 479392 496080 547880 496108
rect 479392 496068 479398 496080
rect 547874 496068 547880 496080
rect 547932 496068 547938 496120
rect 49234 495456 49240 495508
rect 49292 495496 49298 495508
rect 50338 495496 50344 495508
rect 49292 495468 50344 495496
rect 49292 495456 49298 495468
rect 50338 495456 50344 495468
rect 50396 495456 50402 495508
rect 478322 495388 478328 495440
rect 478380 495428 478386 495440
rect 480990 495428 480996 495440
rect 478380 495400 480996 495428
rect 478380 495388 478386 495400
rect 480990 495388 480996 495400
rect 481048 495388 481054 495440
rect 445754 494844 445760 494896
rect 445812 494884 445818 494896
rect 512914 494884 512920 494896
rect 445812 494856 512920 494884
rect 445812 494844 445818 494856
rect 512914 494844 512920 494856
rect 512972 494844 512978 494896
rect 398834 494776 398840 494828
rect 398892 494816 398898 494828
rect 511166 494816 511172 494828
rect 398892 494788 511172 494816
rect 398892 494776 398898 494788
rect 511166 494776 511172 494788
rect 511224 494776 511230 494828
rect 285674 494708 285680 494760
rect 285732 494748 285738 494760
rect 320450 494748 320456 494760
rect 285732 494720 320456 494748
rect 285732 494708 285738 494720
rect 320450 494708 320456 494720
rect 320508 494708 320514 494760
rect 369118 494708 369124 494760
rect 369176 494748 369182 494760
rect 483198 494748 483204 494760
rect 369176 494720 483204 494748
rect 369176 494708 369182 494720
rect 483198 494708 483204 494720
rect 483256 494708 483262 494760
rect 287054 494640 287060 494692
rect 287112 494680 287118 494692
rect 287882 494680 287888 494692
rect 287112 494652 287888 494680
rect 287112 494640 287118 494652
rect 287882 494640 287888 494652
rect 287940 494640 287946 494692
rect 288434 494640 288440 494692
rect 288492 494680 288498 494692
rect 289354 494680 289360 494692
rect 288492 494652 289360 494680
rect 288492 494640 288498 494652
rect 289354 494640 289360 494652
rect 289412 494640 289418 494692
rect 299474 494640 299480 494692
rect 299532 494680 299538 494692
rect 300394 494680 300400 494692
rect 299532 494652 300400 494680
rect 299532 494640 299538 494652
rect 300394 494640 300400 494652
rect 300452 494640 300458 494692
rect 307754 494640 307760 494692
rect 307812 494680 307818 494692
rect 308490 494680 308496 494692
rect 307812 494652 308496 494680
rect 307812 494640 307818 494652
rect 308490 494640 308496 494652
rect 308548 494640 308554 494692
rect 311894 494300 311900 494352
rect 311952 494340 311958 494352
rect 312906 494340 312912 494352
rect 311952 494312 312912 494340
rect 311952 494300 311958 494312
rect 312906 494300 312912 494312
rect 312964 494300 312970 494352
rect 254578 494028 254584 494080
rect 254636 494068 254642 494080
rect 261570 494068 261576 494080
rect 254636 494040 261576 494068
rect 254636 494028 254642 494040
rect 261570 494028 261576 494040
rect 261628 494028 261634 494080
rect 358262 493960 358268 494012
rect 358320 494000 358326 494012
rect 362218 494000 362224 494012
rect 358320 493972 362224 494000
rect 358320 493960 358326 493972
rect 362218 493960 362224 493972
rect 362276 493960 362282 494012
rect 481082 493960 481088 494012
rect 481140 494000 481146 494012
rect 483842 494000 483848 494012
rect 481140 493972 483848 494000
rect 481140 493960 481146 493972
rect 483842 493960 483848 493972
rect 483900 493960 483906 494012
rect 296714 493416 296720 493468
rect 296772 493456 296778 493468
rect 297450 493456 297456 493468
rect 296772 493428 297456 493456
rect 296772 493416 296778 493428
rect 297450 493416 297456 493428
rect 297508 493416 297514 493468
rect 402974 493348 402980 493400
rect 403032 493388 403038 493400
rect 512638 493388 512644 493400
rect 403032 493360 512644 493388
rect 403032 493348 403038 493360
rect 512638 493348 512644 493360
rect 512696 493348 512702 493400
rect 389174 493280 389180 493332
rect 389232 493320 389238 493332
rect 510430 493320 510436 493332
rect 389232 493292 510436 493320
rect 389232 493280 389238 493292
rect 510430 493280 510436 493292
rect 510488 493280 510494 493332
rect 298830 492600 298836 492652
rect 298888 492640 298894 492652
rect 302326 492640 302332 492652
rect 298888 492612 302332 492640
rect 298888 492600 298894 492612
rect 302326 492600 302332 492612
rect 302384 492600 302390 492652
rect 285858 491920 285864 491972
rect 285916 491960 285922 491972
rect 292022 491960 292028 491972
rect 285916 491932 292028 491960
rect 285916 491920 285922 491932
rect 292022 491920 292028 491932
rect 292080 491920 292086 491972
rect 392210 491920 392216 491972
rect 392268 491960 392274 491972
rect 412634 491960 412640 491972
rect 392268 491932 412640 491960
rect 392268 491920 392274 491932
rect 412634 491920 412640 491932
rect 412692 491920 412698 491972
rect 358906 489132 358912 489184
rect 358964 489172 358970 489184
rect 580442 489172 580448 489184
rect 358964 489144 580448 489172
rect 358964 489132 358970 489144
rect 580442 489132 580448 489144
rect 580500 489132 580506 489184
rect 254670 488520 254676 488572
rect 254728 488560 254734 488572
rect 279418 488560 279424 488572
rect 254728 488532 279424 488560
rect 254728 488520 254734 488532
rect 279418 488520 279424 488532
rect 279476 488520 279482 488572
rect 276014 487772 276020 487824
rect 276072 487812 276078 487824
rect 320358 487812 320364 487824
rect 276072 487784 320364 487812
rect 276072 487772 276078 487784
rect 320358 487772 320364 487784
rect 320416 487772 320422 487824
rect 479058 486412 479064 486464
rect 479116 486452 479122 486464
rect 580350 486452 580356 486464
rect 479116 486424 580356 486452
rect 479116 486412 479122 486424
rect 580350 486412 580356 486424
rect 580408 486412 580414 486464
rect 49418 485800 49424 485852
rect 49476 485840 49482 485852
rect 51718 485840 51724 485852
rect 49476 485812 51724 485840
rect 49476 485800 49482 485812
rect 51718 485800 51724 485812
rect 51776 485800 51782 485852
rect 482370 485732 482376 485784
rect 482428 485772 482434 485784
rect 580166 485772 580172 485784
rect 482428 485744 580172 485772
rect 482428 485732 482434 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 364334 482264 364340 482316
rect 364392 482304 364398 482316
rect 497366 482304 497372 482316
rect 364392 482276 497372 482304
rect 364392 482264 364398 482276
rect 497366 482264 497372 482276
rect 497424 482264 497430 482316
rect 254394 481652 254400 481704
rect 254452 481692 254458 481704
rect 268470 481692 268476 481704
rect 254452 481664 268476 481692
rect 254452 481652 254458 481664
rect 268470 481652 268476 481664
rect 268528 481652 268534 481704
rect 49326 481584 49332 481636
rect 49384 481624 49390 481636
rect 50430 481624 50436 481636
rect 49384 481596 50436 481624
rect 49384 481584 49390 481596
rect 50430 481584 50436 481596
rect 50488 481584 50494 481636
rect 310606 480904 310612 480956
rect 310664 480944 310670 480956
rect 350258 480944 350264 480956
rect 310664 480916 350264 480944
rect 310664 480904 310670 480916
rect 350258 480904 350264 480916
rect 350316 480904 350322 480956
rect 382274 480904 382280 480956
rect 382332 480944 382338 480956
rect 506382 480944 506388 480956
rect 382332 480916 506388 480944
rect 382332 480904 382338 480916
rect 506382 480904 506388 480916
rect 506440 480904 506446 480956
rect 373994 479476 374000 479528
rect 374052 479516 374058 479528
rect 471330 479516 471336 479528
rect 374052 479488 471336 479516
rect 374052 479476 374058 479488
rect 471330 479476 471336 479488
rect 471388 479476 471394 479528
rect 385034 478116 385040 478168
rect 385092 478156 385098 478168
rect 460198 478156 460204 478168
rect 385092 478128 460204 478156
rect 385092 478116 385098 478128
rect 460198 478116 460204 478128
rect 460256 478116 460262 478168
rect 391934 476756 391940 476808
rect 391992 476796 391998 476808
rect 480622 476796 480628 476808
rect 391992 476768 480628 476796
rect 391992 476756 391998 476768
rect 480622 476756 480628 476768
rect 480680 476756 480686 476808
rect 254210 476076 254216 476128
rect 254268 476116 254274 476128
rect 265710 476116 265716 476128
rect 254268 476088 265716 476116
rect 254268 476076 254274 476088
rect 265710 476076 265716 476088
rect 265768 476076 265774 476128
rect 46382 473288 46388 473340
rect 46440 473328 46446 473340
rect 48958 473328 48964 473340
rect 46440 473300 48964 473328
rect 46440 473288 46446 473300
rect 48958 473288 48964 473300
rect 49016 473288 49022 473340
rect 338758 471928 338764 471980
rect 338816 471968 338822 471980
rect 580166 471968 580172 471980
rect 338816 471940 580172 471968
rect 338816 471928 338822 471940
rect 580166 471928 580172 471940
rect 580224 471928 580230 471980
rect 254486 470568 254492 470620
rect 254544 470608 254550 470620
rect 264330 470608 264336 470620
rect 254544 470580 264336 470608
rect 254544 470568 254550 470580
rect 264330 470568 264336 470580
rect 264388 470568 264394 470620
rect 45462 467780 45468 467832
rect 45520 467820 45526 467832
rect 48774 467820 48780 467832
rect 45520 467792 48780 467820
rect 45520 467780 45526 467792
rect 48774 467780 48780 467792
rect 48832 467820 48838 467832
rect 49050 467820 49056 467832
rect 48832 467792 49056 467820
rect 48832 467780 48838 467792
rect 49050 467780 49056 467792
rect 49108 467780 49114 467832
rect 254670 465060 254676 465112
rect 254728 465100 254734 465112
rect 289078 465100 289084 465112
rect 254728 465072 289084 465100
rect 254728 465060 254734 465072
rect 289078 465060 289084 465072
rect 289136 465060 289142 465112
rect 47854 462272 47860 462324
rect 47912 462312 47918 462324
rect 50798 462312 50804 462324
rect 47912 462284 50804 462312
rect 47912 462272 47918 462284
rect 50798 462272 50804 462284
rect 50856 462272 50862 462324
rect 297634 460164 297640 460216
rect 297692 460204 297698 460216
rect 313366 460204 313372 460216
rect 297692 460176 313372 460204
rect 297692 460164 297698 460176
rect 313366 460164 313372 460176
rect 313424 460164 313430 460216
rect 254302 458192 254308 458244
rect 254360 458232 254366 458244
rect 269942 458232 269948 458244
rect 254360 458204 269948 458232
rect 254360 458192 254366 458204
rect 269942 458192 269948 458204
rect 270000 458192 270006 458244
rect 46474 456356 46480 456408
rect 46532 456396 46538 456408
rect 49786 456396 49792 456408
rect 46532 456368 49792 456396
rect 46532 456356 46538 456368
rect 49786 456356 49792 456368
rect 49844 456356 49850 456408
rect 299566 453976 299572 454028
rect 299624 454016 299630 454028
rect 300946 454016 300952 454028
rect 299624 453988 300952 454016
rect 299624 453976 299630 453988
rect 300946 453976 300952 453988
rect 301004 453976 301010 454028
rect 254670 452616 254676 452668
rect 254728 452656 254734 452668
rect 284938 452656 284944 452668
rect 254728 452628 284944 452656
rect 254728 452616 254734 452628
rect 284938 452616 284944 452628
rect 284996 452616 285002 452668
rect 50614 450712 50620 450764
rect 50672 450752 50678 450764
rect 51258 450752 51264 450764
rect 50672 450724 51264 450752
rect 50672 450712 50678 450724
rect 51258 450712 51264 450724
rect 51316 450712 51322 450764
rect 254670 447108 254676 447160
rect 254728 447148 254734 447160
rect 278222 447148 278228 447160
rect 254728 447120 278228 447148
rect 254728 447108 254734 447120
rect 278222 447108 278228 447120
rect 278280 447108 278286 447160
rect 46566 445680 46572 445732
rect 46624 445720 46630 445732
rect 48314 445720 48320 445732
rect 46624 445692 48320 445720
rect 46624 445680 46630 445692
rect 48314 445680 48320 445692
rect 48372 445680 48378 445732
rect 254394 441736 254400 441788
rect 254452 441776 254458 441788
rect 257522 441776 257528 441788
rect 254452 441748 257528 441776
rect 254452 441736 254458 441748
rect 257522 441736 257528 441748
rect 257580 441736 257586 441788
rect 46658 438812 46664 438864
rect 46716 438852 46722 438864
rect 48314 438852 48320 438864
rect 46716 438824 48320 438852
rect 46716 438812 46722 438824
rect 48314 438812 48320 438824
rect 48372 438812 48378 438864
rect 254670 434732 254676 434784
rect 254728 434772 254734 434784
rect 291838 434772 291844 434784
rect 254728 434744 291844 434772
rect 254728 434732 254734 434744
rect 291838 434732 291844 434744
rect 291896 434732 291902 434784
rect 46750 433236 46756 433288
rect 46808 433276 46814 433288
rect 49142 433276 49148 433288
rect 46808 433248 49148 433276
rect 46808 433236 46814 433248
rect 49142 433236 49148 433248
rect 49200 433236 49206 433288
rect 518158 431876 518164 431928
rect 518216 431916 518222 431928
rect 579614 431916 579620 431928
rect 518216 431888 579620 431916
rect 518216 431876 518222 431888
rect 579614 431876 579620 431888
rect 579672 431876 579678 431928
rect 254210 429156 254216 429208
rect 254268 429196 254274 429208
rect 351454 429196 351460 429208
rect 254268 429168 351460 429196
rect 254268 429156 254274 429168
rect 351454 429156 351460 429168
rect 351512 429156 351518 429208
rect 46842 427728 46848 427780
rect 46900 427768 46906 427780
rect 49418 427768 49424 427780
rect 46900 427740 49424 427768
rect 46900 427728 46906 427740
rect 49418 427728 49424 427740
rect 49476 427728 49482 427780
rect 254670 423648 254676 423700
rect 254728 423688 254734 423700
rect 323670 423688 323676 423700
rect 254728 423660 323676 423688
rect 254728 423648 254734 423660
rect 323670 423648 323676 423660
rect 323728 423648 323734 423700
rect 323578 419432 323584 419484
rect 323636 419472 323642 419484
rect 580166 419472 580172 419484
rect 323636 419444 580172 419472
rect 323636 419432 323642 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 254394 418140 254400 418192
rect 254452 418180 254458 418192
rect 287698 418180 287704 418192
rect 254452 418152 287704 418180
rect 254452 418140 254458 418152
rect 287698 418140 287704 418152
rect 287756 418140 287762 418192
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 50522 409884 50528 409896
rect 3200 409856 50528 409884
rect 3200 409844 3206 409856
rect 50522 409844 50528 409856
rect 50580 409844 50586 409896
rect 254302 405696 254308 405748
rect 254360 405736 254366 405748
rect 350810 405736 350816 405748
rect 254360 405708 350816 405736
rect 254360 405696 254366 405708
rect 350810 405696 350816 405708
rect 350868 405696 350874 405748
rect 366358 405628 366364 405680
rect 366416 405668 366422 405680
rect 580166 405668 580172 405680
rect 366416 405640 580172 405668
rect 366416 405628 366422 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 254486 400188 254492 400240
rect 254544 400228 254550 400240
rect 350626 400228 350632 400240
rect 254544 400200 350632 400228
rect 254544 400188 254550 400200
rect 350626 400188 350632 400200
rect 350684 400188 350690 400240
rect 254486 394952 254492 395004
rect 254544 394992 254550 395004
rect 260374 394992 260380 395004
rect 254544 394964 260380 394992
rect 254544 394952 254550 394964
rect 260374 394952 260380 394964
rect 260432 394952 260438 395004
rect 46842 391960 46848 392012
rect 46900 392000 46906 392012
rect 48314 392000 48320 392012
rect 46900 391972 48320 392000
rect 46900 391960 46906 391972
rect 48314 391960 48320 391972
rect 48372 391960 48378 392012
rect 254486 389172 254492 389224
rect 254544 389212 254550 389224
rect 313918 389212 313924 389224
rect 254544 389184 313924 389212
rect 254544 389172 254550 389184
rect 313918 389172 313924 389184
rect 313976 389172 313982 389224
rect 46750 385024 46756 385076
rect 46808 385064 46814 385076
rect 48314 385064 48320 385076
rect 46808 385036 48320 385064
rect 46808 385024 46814 385036
rect 48314 385024 48320 385036
rect 48372 385024 48378 385076
rect 254210 382236 254216 382288
rect 254268 382276 254274 382288
rect 289170 382276 289176 382288
rect 254268 382248 289176 382276
rect 254268 382236 254274 382248
rect 289170 382236 289176 382248
rect 289228 382236 289234 382288
rect 46658 379516 46664 379568
rect 46716 379556 46722 379568
rect 49418 379556 49424 379568
rect 46716 379528 49424 379556
rect 46716 379516 46722 379528
rect 49418 379516 49424 379528
rect 49476 379516 49482 379568
rect 254118 376728 254124 376780
rect 254176 376768 254182 376780
rect 350902 376768 350908 376780
rect 254176 376740 350908 376768
rect 254176 376728 254182 376740
rect 350902 376728 350908 376740
rect 350960 376728 350966 376780
rect 254394 371220 254400 371272
rect 254452 371260 254458 371272
rect 301498 371260 301504 371272
rect 254452 371232 301504 371260
rect 254452 371220 254458 371232
rect 301498 371220 301504 371232
rect 301556 371220 301562 371272
rect 254486 365712 254492 365764
rect 254544 365752 254550 365764
rect 287790 365752 287796 365764
rect 254544 365724 287796 365752
rect 254544 365712 254550 365724
rect 287790 365712 287796 365724
rect 287848 365712 287854 365764
rect 320818 365644 320824 365696
rect 320876 365684 320882 365696
rect 580166 365684 580172 365696
rect 320876 365656 580172 365684
rect 320876 365644 320882 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 299658 362176 299664 362228
rect 299716 362216 299722 362228
rect 314654 362216 314660 362228
rect 299716 362188 314660 362216
rect 299716 362176 299722 362188
rect 314654 362176 314660 362188
rect 314712 362176 314718 362228
rect 253934 358844 253940 358896
rect 253992 358884 253998 358896
rect 256142 358884 256148 358896
rect 253992 358856 256148 358884
rect 253992 358844 253998 358856
rect 256142 358844 256148 358856
rect 256200 358844 256206 358896
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 50614 357456 50620 357468
rect 3200 357428 50620 357456
rect 3200 357416 3206 357428
rect 50614 357416 50620 357428
rect 50672 357416 50678 357468
rect 307846 355308 307852 355360
rect 307904 355348 307910 355360
rect 349798 355348 349804 355360
rect 307904 355320 349804 355348
rect 307904 355308 307910 355320
rect 349798 355308 349804 355320
rect 349856 355308 349862 355360
rect 288526 353948 288532 354000
rect 288584 353988 288590 354000
rect 352650 353988 352656 354000
rect 288584 353960 352656 353988
rect 288584 353948 288590 353960
rect 352650 353948 352656 353960
rect 352708 353948 352714 354000
rect 482554 353948 482560 354000
rect 482612 353988 482618 354000
rect 552014 353988 552020 354000
rect 482612 353960 552020 353988
rect 482612 353948 482618 353960
rect 552014 353948 552020 353960
rect 552072 353948 552078 354000
rect 254486 353268 254492 353320
rect 254544 353308 254550 353320
rect 289262 353308 289268 353320
rect 254544 353280 289268 353308
rect 254544 353268 254550 353280
rect 289262 353268 289268 353280
rect 289320 353268 289326 353320
rect 362218 353200 362224 353252
rect 362276 353240 362282 353252
rect 580166 353240 580172 353252
rect 362276 353212 580172 353240
rect 362276 353200 362282 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 498194 352588 498200 352640
rect 498252 352628 498258 352640
rect 510062 352628 510068 352640
rect 498252 352600 510068 352628
rect 498252 352588 498258 352600
rect 510062 352588 510068 352600
rect 510120 352588 510126 352640
rect 287146 352520 287152 352572
rect 287204 352560 287210 352572
rect 350166 352560 350172 352572
rect 287204 352532 350172 352560
rect 287204 352520 287210 352532
rect 350166 352520 350172 352532
rect 350224 352520 350230 352572
rect 431954 352520 431960 352572
rect 432012 352560 432018 352572
rect 512546 352560 512552 352572
rect 432012 352532 512552 352560
rect 432012 352520 432018 352532
rect 512546 352520 512552 352532
rect 512604 352520 512610 352572
rect 289814 351160 289820 351212
rect 289872 351200 289878 351212
rect 319162 351200 319168 351212
rect 289872 351172 319168 351200
rect 289872 351160 289878 351172
rect 319162 351160 319168 351172
rect 319220 351160 319226 351212
rect 258074 349800 258080 349852
rect 258132 349840 258138 349852
rect 511074 349840 511080 349852
rect 258132 349812 511080 349840
rect 258132 349800 258138 349812
rect 511074 349800 511080 349812
rect 511132 349800 511138 349852
rect 299014 348372 299020 348424
rect 299072 348412 299078 348424
rect 307754 348412 307760 348424
rect 299072 348384 307760 348412
rect 299072 348372 299078 348384
rect 307754 348372 307760 348384
rect 307812 348372 307818 348424
rect 254762 347760 254768 347812
rect 254820 347800 254826 347812
rect 346394 347800 346400 347812
rect 254820 347772 346400 347800
rect 254820 347760 254826 347772
rect 346394 347760 346400 347772
rect 346452 347760 346458 347812
rect 288434 347012 288440 347064
rect 288492 347052 288498 347064
rect 352098 347052 352104 347064
rect 288492 347024 352104 347052
rect 288492 347012 288498 347024
rect 352098 347012 352104 347024
rect 352156 347012 352162 347064
rect 282914 345652 282920 345704
rect 282972 345692 282978 345704
rect 319070 345692 319076 345704
rect 282972 345664 319076 345692
rect 282972 345652 282978 345664
rect 319070 345652 319076 345664
rect 319128 345652 319134 345704
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 50246 345080 50252 345092
rect 3384 345052 50252 345080
rect 3384 345040 3390 345052
rect 50246 345040 50252 345052
rect 50304 345040 50310 345092
rect 297818 344360 297824 344412
rect 297876 344400 297882 344412
rect 311986 344400 311992 344412
rect 297876 344372 311992 344400
rect 297876 344360 297882 344372
rect 311986 344360 311992 344372
rect 312044 344360 312050 344412
rect 271874 344292 271880 344344
rect 271932 344332 271938 344344
rect 318978 344332 318984 344344
rect 271932 344304 318984 344332
rect 271932 344292 271938 344304
rect 318978 344292 318984 344304
rect 319036 344292 319042 344344
rect 283098 342864 283104 342916
rect 283156 342904 283162 342916
rect 349890 342904 349896 342916
rect 283156 342876 349896 342904
rect 283156 342864 283162 342876
rect 349890 342864 349896 342876
rect 349948 342864 349954 342916
rect 254670 342252 254676 342304
rect 254728 342292 254734 342304
rect 296162 342292 296168 342304
rect 254728 342264 296168 342292
rect 254728 342252 254734 342264
rect 296162 342252 296168 342264
rect 296220 342252 296226 342304
rect 296806 341640 296812 341692
rect 296864 341680 296870 341692
rect 311986 341680 311992 341692
rect 296864 341652 311992 341680
rect 296864 341640 296870 341652
rect 311986 341640 311992 341652
rect 312044 341640 312050 341692
rect 303798 341572 303804 341624
rect 303856 341612 303862 341624
rect 320266 341612 320272 341624
rect 303856 341584 320272 341612
rect 303856 341572 303862 341584
rect 320266 341572 320272 341584
rect 320324 341572 320330 341624
rect 285766 341504 285772 341556
rect 285824 341544 285830 341556
rect 352466 341544 352472 341556
rect 285824 341516 352472 341544
rect 285824 341504 285830 341516
rect 352466 341504 352472 341516
rect 352524 341504 352530 341556
rect 478966 341504 478972 341556
rect 479024 341544 479030 341556
rect 580350 341544 580356 341556
rect 479024 341516 580356 341544
rect 479024 341504 479030 341516
rect 580350 341504 580356 341516
rect 580408 341504 580414 341556
rect 296714 340144 296720 340196
rect 296772 340184 296778 340196
rect 349706 340184 349712 340196
rect 296772 340156 349712 340184
rect 296772 340144 296778 340156
rect 349706 340144 349712 340156
rect 349764 340144 349770 340196
rect 267734 338784 267740 338836
rect 267792 338824 267798 338836
rect 318886 338824 318892 338836
rect 267792 338796 318892 338824
rect 267792 338784 267798 338796
rect 318886 338784 318892 338796
rect 318944 338784 318950 338836
rect 289906 338716 289912 338768
rect 289964 338756 289970 338768
rect 352282 338756 352288 338768
rect 289964 338728 352288 338756
rect 289964 338716 289970 338728
rect 352282 338716 352288 338728
rect 352340 338716 352346 338768
rect 299474 337492 299480 337544
rect 299532 337532 299538 337544
rect 319346 337532 319352 337544
rect 299532 337504 319352 337532
rect 299532 337492 299538 337504
rect 319346 337492 319352 337504
rect 319404 337492 319410 337544
rect 260834 337356 260840 337408
rect 260892 337396 260898 337408
rect 319254 337396 319260 337408
rect 260892 337368 319260 337396
rect 260892 337356 260898 337368
rect 319254 337356 319260 337368
rect 319312 337356 319318 337408
rect 254762 335996 254768 336048
rect 254820 336036 254826 336048
rect 350718 336036 350724 336048
rect 254820 336008 350724 336036
rect 254820 335996 254826 336008
rect 350718 335996 350724 336008
rect 350776 335996 350782 336048
rect 313918 335384 313924 335436
rect 313976 335424 313982 335436
rect 318058 335424 318064 335436
rect 313976 335396 318064 335424
rect 313976 335384 313982 335396
rect 318058 335384 318064 335396
rect 318116 335384 318122 335436
rect 254670 335316 254676 335368
rect 254728 335356 254734 335368
rect 332226 335356 332232 335368
rect 254728 335328 332232 335356
rect 254728 335316 254734 335328
rect 332226 335316 332232 335328
rect 332284 335316 332290 335368
rect 298554 334704 298560 334756
rect 298612 334744 298618 334756
rect 311894 334744 311900 334756
rect 298612 334716 311900 334744
rect 298612 334704 298618 334716
rect 311894 334704 311900 334716
rect 311952 334704 311958 334756
rect 310514 334636 310520 334688
rect 310572 334676 310578 334688
rect 352006 334676 352012 334688
rect 310572 334648 352012 334676
rect 310572 334636 310578 334648
rect 352006 334636 352012 334648
rect 352064 334636 352070 334688
rect 291286 334568 291292 334620
rect 291344 334608 291350 334620
rect 351086 334608 351092 334620
rect 291344 334580 351092 334608
rect 291344 334568 291350 334580
rect 351086 334568 351092 334580
rect 351144 334568 351150 334620
rect 306466 333344 306472 333396
rect 306524 333384 306530 333396
rect 350994 333384 351000 333396
rect 306524 333356 351000 333384
rect 306524 333344 306530 333356
rect 350994 333344 351000 333356
rect 351052 333344 351058 333396
rect 286318 333276 286324 333328
rect 286376 333316 286382 333328
rect 352374 333316 352380 333328
rect 286376 333288 352380 333316
rect 286376 333276 286382 333288
rect 352374 333276 352380 333288
rect 352432 333276 352438 333328
rect 298002 333208 298008 333260
rect 298060 333248 298066 333260
rect 320174 333248 320180 333260
rect 298060 333220 320180 333248
rect 298060 333208 298066 333220
rect 320174 333208 320180 333220
rect 320232 333208 320238 333260
rect 301498 333140 301504 333192
rect 301556 333180 301562 333192
rect 306466 333180 306472 333192
rect 301556 333152 306472 333180
rect 301556 333140 301562 333152
rect 306466 333140 306472 333152
rect 306524 333140 306530 333192
rect 285122 332188 285128 332240
rect 285180 332228 285186 332240
rect 323210 332228 323216 332240
rect 285180 332200 323216 332228
rect 285180 332188 285186 332200
rect 323210 332188 323216 332200
rect 323268 332188 323274 332240
rect 296438 332120 296444 332172
rect 296496 332160 296502 332172
rect 305086 332160 305092 332172
rect 296496 332132 305092 332160
rect 296496 332120 296502 332132
rect 305086 332120 305092 332132
rect 305144 332120 305150 332172
rect 349706 332120 349712 332172
rect 349764 332160 349770 332172
rect 349982 332160 349988 332172
rect 349764 332132 349988 332160
rect 349764 332120 349770 332132
rect 349982 332120 349988 332132
rect 350040 332120 350046 332172
rect 295150 332052 295156 332104
rect 295208 332092 295214 332104
rect 306374 332092 306380 332104
rect 295208 332064 306380 332092
rect 295208 332052 295214 332064
rect 306374 332052 306380 332064
rect 306432 332052 306438 332104
rect 296346 331984 296352 332036
rect 296404 332024 296410 332036
rect 309134 332024 309140 332036
rect 296404 331996 309140 332024
rect 296404 331984 296410 331996
rect 309134 331984 309140 331996
rect 309192 331984 309198 332036
rect 294966 331916 294972 331968
rect 295024 331956 295030 331968
rect 309226 331956 309232 331968
rect 295024 331928 309232 331956
rect 295024 331916 295030 331928
rect 309226 331916 309232 331928
rect 309284 331916 309290 331968
rect 295058 331848 295064 331900
rect 295116 331888 295122 331900
rect 302418 331888 302424 331900
rect 295116 331860 302424 331888
rect 295116 331848 295122 331860
rect 302418 331848 302424 331860
rect 302476 331848 302482 331900
rect 303614 331848 303620 331900
rect 303672 331888 303678 331900
rect 350350 331888 350356 331900
rect 303672 331860 350356 331888
rect 303672 331848 303678 331860
rect 350350 331848 350356 331860
rect 350408 331848 350414 331900
rect 323670 331780 323676 331832
rect 323728 331820 323734 331832
rect 325142 331820 325148 331832
rect 323728 331792 325148 331820
rect 323728 331780 323734 331792
rect 325142 331780 325148 331792
rect 325200 331780 325206 331832
rect 293862 331712 293868 331764
rect 293920 331752 293926 331764
rect 309042 331752 309048 331764
rect 293920 331724 309048 331752
rect 293920 331712 293926 331724
rect 309042 331712 309048 331724
rect 309100 331712 309106 331764
rect 298738 331644 298744 331696
rect 298796 331684 298802 331696
rect 343818 331684 343824 331696
rect 298796 331656 343824 331684
rect 298796 331644 298802 331656
rect 343818 331644 343824 331656
rect 343876 331644 343882 331696
rect 296254 331576 296260 331628
rect 296312 331616 296318 331628
rect 313550 331616 313556 331628
rect 296312 331588 313556 331616
rect 296312 331576 296318 331588
rect 313550 331576 313556 331588
rect 313608 331576 313614 331628
rect 292114 331508 292120 331560
rect 292172 331548 292178 331560
rect 321922 331548 321928 331560
rect 292172 331520 321928 331548
rect 292172 331508 292178 331520
rect 321922 331508 321928 331520
rect 321980 331508 321986 331560
rect 327718 331508 327724 331560
rect 327776 331548 327782 331560
rect 333514 331548 333520 331560
rect 327776 331520 333520 331548
rect 327776 331508 327782 331520
rect 333514 331508 333520 331520
rect 333572 331508 333578 331560
rect 338022 331508 338028 331560
rect 338080 331548 338086 331560
rect 353570 331548 353576 331560
rect 338080 331520 353576 331548
rect 338080 331508 338086 331520
rect 353570 331508 353576 331520
rect 353628 331508 353634 331560
rect 298830 331440 298836 331492
rect 298888 331480 298894 331492
rect 329006 331480 329012 331492
rect 298888 331452 329012 331480
rect 298888 331440 298894 331452
rect 329006 331440 329012 331452
rect 329064 331440 329070 331492
rect 339310 331440 339316 331492
rect 339368 331480 339374 331492
rect 352190 331480 352196 331492
rect 339368 331452 352196 331480
rect 339368 331440 339374 331452
rect 352190 331440 352196 331452
rect 352248 331440 352254 331492
rect 293770 331372 293776 331424
rect 293828 331412 293834 331424
rect 330938 331412 330944 331424
rect 293828 331384 330944 331412
rect 293828 331372 293834 331384
rect 330938 331372 330944 331384
rect 330996 331372 331002 331424
rect 336090 331372 336096 331424
rect 336148 331412 336154 331424
rect 354674 331412 354680 331424
rect 336148 331384 354680 331412
rect 336148 331372 336154 331384
rect 354674 331372 354680 331384
rect 354732 331372 354738 331424
rect 298922 331304 298928 331356
rect 298980 331344 298986 331356
rect 307754 331344 307760 331356
rect 298980 331316 307760 331344
rect 298980 331304 298986 331316
rect 307754 331304 307760 331316
rect 307812 331304 307818 331356
rect 327718 331304 327724 331356
rect 327776 331344 327782 331356
rect 353662 331344 353668 331356
rect 327776 331316 353668 331344
rect 327776 331304 327782 331316
rect 353662 331304 353668 331316
rect 353720 331304 353726 331356
rect 293678 331236 293684 331288
rect 293736 331276 293742 331288
rect 301958 331276 301964 331288
rect 293736 331248 301964 331276
rect 293736 331236 293742 331248
rect 301958 331236 301964 331248
rect 302016 331236 302022 331288
rect 345106 331236 345112 331288
rect 345164 331276 345170 331288
rect 354766 331276 354772 331288
rect 345164 331248 354772 331276
rect 345164 331236 345170 331248
rect 354766 331236 354772 331248
rect 354824 331236 354830 331288
rect 284294 330488 284300 330540
rect 284352 330528 284358 330540
rect 286318 330528 286324 330540
rect 284352 330500 286324 330528
rect 284352 330488 284358 330500
rect 286318 330488 286324 330500
rect 286376 330488 286382 330540
rect 299198 330080 299204 330132
rect 299256 330120 299262 330132
rect 326430 330120 326436 330132
rect 299256 330092 326436 330120
rect 299256 330080 299262 330092
rect 326430 330080 326436 330092
rect 326488 330080 326494 330132
rect 299290 330012 299296 330064
rect 299348 330052 299354 330064
rect 334526 330052 334532 330064
rect 299348 330024 334532 330052
rect 299348 330012 299354 330024
rect 334526 330012 334532 330024
rect 334584 330012 334590 330064
rect 299106 329944 299112 329996
rect 299164 329984 299170 329996
rect 340230 329984 340236 329996
rect 299164 329956 340236 329984
rect 299164 329944 299170 329956
rect 340230 329944 340236 329956
rect 340288 329944 340294 329996
rect 254210 329876 254216 329928
rect 254268 329916 254274 329928
rect 285030 329916 285036 329928
rect 254268 329888 285036 329916
rect 254268 329876 254274 329888
rect 285030 329876 285036 329888
rect 285088 329876 285094 329928
rect 299382 329876 299388 329928
rect 299440 329916 299446 329928
rect 347406 329916 347412 329928
rect 299440 329888 347412 329916
rect 299440 329876 299446 329888
rect 347406 329876 347412 329888
rect 347464 329876 347470 329928
rect 254670 329808 254676 329860
rect 254728 329848 254734 329860
rect 350074 329848 350080 329860
rect 254728 329820 350080 329848
rect 254728 329808 254734 329820
rect 350074 329808 350080 329820
rect 350132 329808 350138 329860
rect 254486 325592 254492 325644
rect 254544 325632 254550 325644
rect 292114 325632 292120 325644
rect 254544 325604 292120 325632
rect 254544 325592 254550 325604
rect 292114 325592 292120 325604
rect 292172 325592 292178 325644
rect 349798 325048 349804 325100
rect 349856 325048 349862 325100
rect 349890 325048 349896 325100
rect 349948 325048 349954 325100
rect 349816 324896 349844 325048
rect 349908 324896 349936 325048
rect 349798 324844 349804 324896
rect 349856 324844 349862 324896
rect 349890 324844 349896 324896
rect 349948 324844 349954 324896
rect 281534 324232 281540 324284
rect 281592 324272 281598 324284
rect 297726 324272 297732 324284
rect 281592 324244 297732 324272
rect 281592 324232 281598 324244
rect 297726 324232 297732 324244
rect 297784 324232 297790 324284
rect 254302 320084 254308 320136
rect 254360 320124 254366 320136
rect 285122 320124 285128 320136
rect 254360 320096 285128 320124
rect 254360 320084 254366 320096
rect 285122 320084 285128 320096
rect 285180 320084 285186 320136
rect 287790 318724 287796 318776
rect 287848 318764 287854 318776
rect 297726 318764 297732 318776
rect 287848 318736 297732 318764
rect 287848 318724 287854 318736
rect 297726 318724 297732 318736
rect 297784 318724 297790 318776
rect 285030 317364 285036 317416
rect 285088 317404 285094 317416
rect 297726 317404 297732 317416
rect 285088 317376 297732 317404
rect 285088 317364 285094 317376
rect 297726 317364 297732 317376
rect 297784 317364 297790 317416
rect 297266 316004 297272 316056
rect 297324 316044 297330 316056
rect 297726 316044 297732 316056
rect 297324 316016 297732 316044
rect 297324 316004 297330 316016
rect 297726 316004 297732 316016
rect 297784 316004 297790 316056
rect 351362 314644 351368 314696
rect 351420 314684 351426 314696
rect 351914 314684 351920 314696
rect 351420 314656 351920 314684
rect 351420 314644 351426 314656
rect 351914 314644 351920 314656
rect 351972 314644 351978 314696
rect 292850 313216 292856 313268
rect 292908 313256 292914 313268
rect 297910 313256 297916 313268
rect 292908 313228 297916 313256
rect 292908 313216 292914 313228
rect 297910 313216 297916 313228
rect 297968 313216 297974 313268
rect 354030 313216 354036 313268
rect 354088 313256 354094 313268
rect 580166 313256 580172 313268
rect 354088 313228 580172 313256
rect 354088 313216 354094 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 260374 307708 260380 307760
rect 260432 307748 260438 307760
rect 298002 307748 298008 307760
rect 260432 307720 298008 307748
rect 260432 307708 260438 307720
rect 298002 307708 298008 307720
rect 298060 307708 298066 307760
rect 254210 306348 254216 306400
rect 254268 306388 254274 306400
rect 293310 306388 293316 306400
rect 254268 306360 293316 306388
rect 254268 306348 254274 306360
rect 293310 306348 293316 306360
rect 293368 306348 293374 306400
rect 256142 306280 256148 306332
rect 256200 306320 256206 306332
rect 298002 306320 298008 306332
rect 256200 306292 298008 306320
rect 256200 306280 256206 306292
rect 298002 306280 298008 306292
rect 298060 306280 298066 306332
rect 349982 303628 349988 303680
rect 350040 303668 350046 303680
rect 351914 303668 351920 303680
rect 350040 303640 351920 303668
rect 350040 303628 350046 303640
rect 351914 303628 351920 303640
rect 351972 303628 351978 303680
rect 293954 303492 293960 303544
rect 294012 303532 294018 303544
rect 298002 303532 298008 303544
rect 294012 303504 298008 303532
rect 294012 303492 294018 303504
rect 298002 303492 298008 303504
rect 298060 303492 298066 303544
rect 292574 303152 292580 303204
rect 292632 303192 292638 303204
rect 294690 303192 294696 303204
rect 292632 303164 294696 303192
rect 292632 303152 292638 303164
rect 294690 303152 294696 303164
rect 294748 303152 294754 303204
rect 254670 300840 254676 300892
rect 254728 300880 254734 300892
rect 294782 300880 294788 300892
rect 254728 300852 294788 300880
rect 254728 300840 254734 300852
rect 294782 300840 294788 300852
rect 294840 300840 294846 300892
rect 383194 299412 383200 299464
rect 383252 299452 383258 299464
rect 579614 299452 579620 299464
rect 383252 299424 579620 299452
rect 383252 299412 383258 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 254670 295332 254676 295384
rect 254728 295372 254734 295384
rect 285030 295372 285036 295384
rect 254728 295344 285036 295372
rect 254728 295332 254734 295344
rect 285030 295332 285036 295344
rect 285088 295332 285094 295384
rect 297818 295128 297824 295180
rect 297876 295168 297882 295180
rect 299750 295168 299756 295180
rect 297876 295140 299756 295168
rect 297876 295128 297882 295140
rect 299750 295128 299756 295140
rect 299808 295128 299814 295180
rect 286318 292476 286324 292528
rect 286376 292516 286382 292528
rect 298002 292516 298008 292528
rect 286376 292488 298008 292516
rect 286376 292476 286382 292488
rect 298002 292476 298008 292488
rect 298060 292476 298066 292528
rect 295426 289620 295432 289672
rect 295484 289660 295490 289672
rect 298002 289660 298008 289672
rect 295484 289632 298008 289660
rect 295484 289620 295490 289632
rect 298002 289620 298008 289632
rect 298060 289620 298066 289672
rect 292022 288328 292028 288380
rect 292080 288368 292086 288380
rect 298002 288368 298008 288380
rect 292080 288340 298008 288368
rect 292080 288328 292086 288340
rect 298002 288328 298008 288340
rect 298060 288328 298066 288380
rect 297818 287376 297824 287428
rect 297876 287376 297882 287428
rect 297836 287088 297864 287376
rect 297818 287036 297824 287088
rect 297876 287036 297882 287088
rect 297818 285880 297824 285932
rect 297876 285880 297882 285932
rect 297836 285728 297864 285880
rect 297818 285676 297824 285728
rect 297876 285676 297882 285728
rect 289170 285608 289176 285660
rect 289228 285648 289234 285660
rect 297910 285648 297916 285660
rect 289228 285620 297916 285648
rect 289228 285608 289234 285620
rect 297910 285608 297916 285620
rect 297968 285608 297974 285660
rect 254302 282888 254308 282940
rect 254360 282928 254366 282940
rect 264422 282928 264428 282940
rect 254360 282900 264428 282928
rect 254360 282888 254366 282900
rect 264422 282888 264428 282900
rect 264480 282888 264486 282940
rect 3510 282004 3516 282056
rect 3568 282044 3574 282056
rect 295426 282044 295432 282056
rect 3568 282016 295432 282044
rect 3568 282004 3574 282016
rect 295426 282004 295432 282016
rect 295484 282004 295490 282056
rect 50614 281936 50620 281988
rect 50672 281976 50678 281988
rect 296070 281976 296076 281988
rect 50672 281948 296076 281976
rect 50672 281936 50678 281948
rect 296070 281936 296076 281948
rect 296128 281936 296134 281988
rect 46750 281868 46756 281920
rect 46808 281908 46814 281920
rect 279878 281908 279884 281920
rect 46808 281880 279884 281908
rect 46808 281868 46814 281880
rect 279878 281868 279884 281880
rect 279936 281868 279942 281920
rect 48774 281800 48780 281852
rect 48832 281840 48838 281852
rect 52914 281840 52920 281852
rect 48832 281812 52920 281840
rect 48832 281800 48838 281812
rect 52914 281800 52920 281812
rect 52972 281800 52978 281852
rect 3418 281460 3424 281512
rect 3476 281500 3482 281512
rect 500586 281500 500592 281512
rect 3476 281472 500592 281500
rect 3476 281460 3482 281472
rect 500586 281460 500592 281472
rect 500644 281460 500650 281512
rect 50522 281392 50528 281444
rect 50580 281432 50586 281444
rect 512454 281432 512460 281444
rect 50580 281404 512460 281432
rect 50580 281392 50586 281404
rect 512454 281392 512460 281404
rect 512512 281392 512518 281444
rect 49142 281324 49148 281376
rect 49200 281364 49206 281376
rect 281166 281364 281172 281376
rect 49200 281336 281172 281364
rect 49200 281324 49206 281336
rect 281166 281324 281172 281336
rect 281224 281324 281230 281376
rect 285030 281324 285036 281376
rect 285088 281364 285094 281376
rect 352006 281364 352012 281376
rect 285088 281336 352012 281364
rect 285088 281324 285094 281336
rect 352006 281324 352012 281336
rect 352064 281324 352070 281376
rect 48958 281256 48964 281308
rect 49016 281296 49022 281308
rect 51902 281296 51908 281308
rect 49016 281268 51908 281296
rect 49016 281256 49022 281268
rect 51902 281256 51908 281268
rect 51960 281256 51966 281308
rect 54478 281296 54484 281308
rect 52012 281268 54484 281296
rect 49050 281120 49056 281172
rect 49108 281160 49114 281172
rect 52012 281160 52040 281268
rect 54478 281256 54484 281268
rect 54536 281256 54542 281308
rect 55858 281256 55864 281308
rect 55916 281296 55922 281308
rect 279786 281296 279792 281308
rect 55916 281268 279792 281296
rect 55916 281256 55922 281268
rect 279786 281256 279792 281268
rect 279844 281256 279850 281308
rect 52086 281188 52092 281240
rect 52144 281228 52150 281240
rect 280982 281228 280988 281240
rect 52144 281200 280988 281228
rect 52144 281188 52150 281200
rect 280982 281188 280988 281200
rect 281040 281188 281046 281240
rect 280798 281160 280804 281172
rect 49108 281132 52040 281160
rect 52472 281132 280804 281160
rect 49108 281120 49114 281132
rect 48682 281052 48688 281104
rect 48740 281092 48746 281104
rect 52472 281092 52500 281132
rect 280798 281120 280804 281132
rect 280856 281120 280862 281172
rect 48740 281064 52500 281092
rect 48740 281052 48746 281064
rect 52914 281052 52920 281104
rect 52972 281092 52978 281104
rect 278314 281092 278320 281104
rect 52972 281064 278320 281092
rect 52972 281052 52978 281064
rect 278314 281052 278320 281064
rect 278372 281052 278378 281104
rect 49234 280984 49240 281036
rect 49292 281024 49298 281036
rect 276658 281024 276664 281036
rect 49292 280996 55996 281024
rect 49292 280984 49298 280996
rect 48038 280916 48044 280968
rect 48096 280956 48102 280968
rect 55858 280956 55864 280968
rect 48096 280928 55864 280956
rect 48096 280916 48102 280928
rect 55858 280916 55864 280928
rect 55916 280916 55922 280968
rect 55968 280956 55996 280996
rect 57946 280996 276664 281024
rect 57946 280956 57974 280996
rect 276658 280984 276664 280996
rect 276716 280984 276722 281036
rect 55968 280928 57974 280956
rect 254026 280916 254032 280968
rect 254084 280956 254090 280968
rect 351454 280956 351460 280968
rect 254084 280928 351460 280956
rect 254084 280916 254090 280928
rect 351454 280916 351460 280928
rect 351512 280916 351518 280968
rect 51902 280780 51908 280832
rect 51960 280820 51966 280832
rect 53098 280820 53104 280832
rect 51960 280792 53104 280820
rect 51960 280780 51966 280792
rect 53098 280780 53104 280792
rect 53156 280780 53162 280832
rect 297726 280576 297732 280628
rect 297784 280616 297790 280628
rect 300118 280616 300124 280628
rect 297784 280588 300124 280616
rect 297784 280576 297790 280588
rect 300118 280576 300124 280588
rect 300176 280576 300182 280628
rect 347314 280576 347320 280628
rect 347372 280616 347378 280628
rect 350074 280616 350080 280628
rect 347372 280588 350080 280616
rect 347372 280576 347378 280588
rect 350074 280576 350080 280588
rect 350132 280576 350138 280628
rect 50246 280100 50252 280152
rect 50304 280140 50310 280152
rect 478138 280140 478144 280152
rect 50304 280112 478144 280140
rect 50304 280100 50310 280112
rect 478138 280100 478144 280112
rect 478196 280100 478202 280152
rect 3602 280032 3608 280084
rect 3660 280072 3666 280084
rect 405090 280072 405096 280084
rect 3660 280044 405096 280072
rect 3660 280032 3666 280044
rect 405090 280032 405096 280044
rect 405148 280032 405154 280084
rect 46658 279964 46664 280016
rect 46716 280004 46722 280016
rect 279694 280004 279700 280016
rect 46716 279976 279700 280004
rect 46716 279964 46722 279976
rect 279694 279964 279700 279976
rect 279752 279964 279758 280016
rect 299842 279964 299848 280016
rect 299900 280004 299906 280016
rect 304994 280004 305000 280016
rect 299900 279976 305000 280004
rect 299900 279964 299906 279976
rect 304994 279964 305000 279976
rect 305052 279964 305058 280016
rect 46842 279896 46848 279948
rect 46900 279936 46906 279948
rect 279510 279936 279516 279948
rect 46900 279908 279516 279936
rect 46900 279896 46906 279908
rect 279510 279896 279516 279908
rect 279568 279896 279574 279948
rect 298922 279896 298928 279948
rect 298980 279936 298986 279948
rect 303798 279936 303804 279948
rect 298980 279908 303804 279936
rect 298980 279896 298986 279908
rect 303798 279896 303804 279908
rect 303856 279896 303862 279948
rect 48222 279828 48228 279880
rect 48280 279868 48286 279880
rect 279602 279868 279608 279880
rect 48280 279840 279608 279868
rect 48280 279828 48286 279840
rect 279602 279828 279608 279840
rect 279660 279828 279666 279880
rect 296254 279488 296260 279540
rect 296312 279528 296318 279540
rect 310514 279528 310520 279540
rect 296312 279500 310520 279528
rect 296312 279488 296318 279500
rect 310514 279488 310520 279500
rect 310572 279488 310578 279540
rect 59538 279420 59544 279472
rect 59596 279460 59602 279472
rect 297358 279460 297364 279472
rect 59596 279432 297364 279460
rect 59596 279420 59602 279432
rect 297358 279420 297364 279432
rect 297416 279420 297422 279472
rect 321646 279420 321652 279472
rect 321704 279460 321710 279472
rect 352190 279460 352196 279472
rect 321704 279432 352196 279460
rect 321704 279420 321710 279432
rect 352190 279420 352196 279432
rect 352248 279420 352254 279472
rect 289262 279012 289268 279064
rect 289320 279052 289326 279064
rect 315482 279052 315488 279064
rect 289320 279024 315488 279052
rect 289320 279012 289326 279024
rect 315482 279012 315488 279024
rect 315540 279012 315546 279064
rect 287698 278944 287704 278996
rect 287756 278984 287762 278996
rect 321278 278984 321284 278996
rect 287756 278956 321284 278984
rect 287756 278944 287762 278956
rect 321278 278944 321284 278956
rect 321336 278944 321342 278996
rect 296162 278876 296168 278928
rect 296220 278916 296226 278928
rect 330938 278916 330944 278928
rect 296220 278888 330944 278916
rect 296220 278876 296226 278888
rect 330938 278876 330944 278888
rect 330996 278876 331002 278928
rect 294782 278808 294788 278860
rect 294840 278848 294846 278860
rect 342530 278848 342536 278860
rect 294840 278820 342536 278848
rect 294840 278808 294846 278820
rect 342530 278808 342536 278820
rect 342588 278808 342594 278860
rect 293310 278740 293316 278792
rect 293368 278780 293374 278792
rect 349614 278780 349620 278792
rect 293368 278752 349620 278780
rect 293368 278740 293374 278752
rect 349614 278740 349620 278752
rect 349672 278740 349678 278792
rect 295058 278672 295064 278724
rect 295116 278712 295122 278724
rect 345750 278712 345756 278724
rect 295116 278684 345756 278712
rect 295116 278672 295122 278684
rect 345750 278672 345756 278684
rect 345808 278672 345814 278724
rect 296346 278604 296352 278656
rect 296404 278644 296410 278656
rect 296404 278616 337332 278644
rect 296404 278604 296410 278616
rect 296438 278536 296444 278588
rect 296496 278576 296502 278588
rect 296496 278548 336688 278576
rect 296496 278536 296502 278548
rect 295334 278468 295340 278520
rect 295392 278508 295398 278520
rect 335446 278508 335452 278520
rect 295392 278480 335452 278508
rect 295392 278468 295398 278480
rect 335446 278468 335452 278480
rect 335504 278468 335510 278520
rect 294966 278400 294972 278452
rect 295024 278440 295030 278452
rect 322566 278440 322572 278452
rect 295024 278412 322572 278440
rect 295024 278400 295030 278412
rect 322566 278400 322572 278412
rect 322624 278400 322630 278452
rect 336660 278440 336688 278548
rect 337304 278508 337332 278616
rect 337378 278604 337384 278656
rect 337436 278644 337442 278656
rect 341242 278644 341248 278656
rect 337436 278616 341248 278644
rect 337436 278604 337442 278616
rect 341242 278604 341248 278616
rect 341300 278604 341306 278656
rect 339954 278508 339960 278520
rect 337304 278480 339960 278508
rect 339954 278468 339960 278480
rect 340012 278468 340018 278520
rect 338022 278440 338028 278452
rect 336660 278412 338028 278440
rect 338022 278400 338028 278412
rect 338080 278400 338086 278452
rect 294690 278332 294696 278384
rect 294748 278372 294754 278384
rect 319990 278372 319996 278384
rect 294748 278344 319996 278372
rect 294748 278332 294754 278344
rect 319990 278332 319996 278344
rect 320048 278332 320054 278384
rect 295150 278264 295156 278316
rect 295208 278304 295214 278316
rect 318058 278304 318064 278316
rect 295208 278276 318064 278304
rect 295208 278264 295214 278276
rect 318058 278264 318064 278276
rect 318116 278264 318122 278316
rect 287054 278196 287060 278248
rect 287112 278236 287118 278248
rect 287112 278208 299888 278236
rect 287112 278196 287118 278208
rect 295978 278128 295984 278180
rect 296036 278168 296042 278180
rect 296036 278140 296714 278168
rect 296036 278128 296042 278140
rect 296686 277964 296714 278140
rect 299860 278100 299888 278208
rect 300026 278196 300032 278248
rect 300084 278236 300090 278248
rect 305638 278236 305644 278248
rect 300084 278208 305644 278236
rect 300084 278196 300090 278208
rect 305638 278196 305644 278208
rect 305696 278196 305702 278248
rect 303890 278100 303896 278112
rect 299860 278072 303896 278100
rect 303890 278060 303896 278072
rect 303948 278060 303954 278112
rect 334158 278060 334164 278112
rect 334216 278100 334222 278112
rect 338206 278100 338212 278112
rect 334216 278072 338212 278100
rect 334216 278060 334222 278072
rect 338206 278060 338212 278072
rect 338264 278060 338270 278112
rect 341518 278060 341524 278112
rect 341576 278100 341582 278112
rect 351914 278100 351920 278112
rect 341576 278072 351920 278100
rect 341576 278060 341582 278072
rect 351914 278060 351920 278072
rect 351972 278060 351978 278112
rect 298646 277992 298652 278044
rect 298704 278032 298710 278044
rect 303706 278032 303712 278044
rect 298704 278004 303712 278032
rect 298704 277992 298710 278004
rect 303706 277992 303712 278004
rect 303764 277992 303770 278044
rect 317414 277992 317420 278044
rect 317472 278032 317478 278044
rect 343818 278032 343824 278044
rect 317472 278004 343824 278032
rect 317472 277992 317478 278004
rect 343818 277992 343824 278004
rect 343876 277992 343882 278044
rect 301314 277964 301320 277976
rect 296686 277936 301320 277964
rect 301314 277924 301320 277936
rect 301372 277924 301378 277976
rect 308398 277924 308404 277976
rect 308456 277964 308462 277976
rect 313274 277964 313280 277976
rect 308456 277936 313280 277964
rect 308456 277924 308462 277936
rect 313274 277924 313280 277936
rect 313332 277924 313338 277976
rect 316770 277924 316776 277976
rect 316828 277964 316834 277976
rect 323118 277964 323124 277976
rect 316828 277936 323124 277964
rect 316828 277924 316834 277936
rect 323118 277924 323124 277936
rect 323176 277924 323182 277976
rect 323854 277516 323860 277568
rect 323912 277556 323918 277568
rect 326338 277556 326344 277568
rect 323912 277528 326344 277556
rect 323912 277516 323918 277528
rect 326338 277516 326344 277528
rect 326396 277516 326402 277568
rect 324314 277380 324320 277432
rect 324372 277420 324378 277432
rect 327074 277420 327080 277432
rect 324372 277392 327080 277420
rect 324372 277380 324378 277392
rect 327074 277380 327080 277392
rect 327132 277380 327138 277432
rect 297450 276700 297456 276752
rect 297508 276740 297514 276752
rect 309134 276740 309140 276752
rect 297508 276712 309140 276740
rect 297508 276700 297514 276712
rect 309134 276700 309140 276712
rect 309192 276700 309198 276752
rect 314746 276700 314752 276752
rect 314804 276740 314810 276752
rect 350902 276740 350908 276752
rect 314804 276712 350908 276740
rect 314804 276700 314810 276712
rect 350902 276700 350908 276712
rect 350960 276700 350966 276752
rect 8938 276632 8944 276684
rect 8996 276672 9002 276684
rect 485774 276672 485780 276684
rect 8996 276644 485780 276672
rect 8996 276632 9002 276644
rect 485774 276632 485780 276644
rect 485832 276632 485838 276684
rect 297910 276020 297916 276072
rect 297968 276060 297974 276072
rect 298830 276060 298836 276072
rect 297968 276032 298836 276060
rect 297968 276020 297974 276032
rect 298830 276020 298836 276032
rect 298888 276020 298894 276072
rect 297174 275340 297180 275392
rect 297232 275380 297238 275392
rect 311158 275380 311164 275392
rect 297232 275352 311164 275380
rect 297232 275340 297238 275352
rect 311158 275340 311164 275352
rect 311216 275340 311222 275392
rect 299566 275272 299572 275324
rect 299624 275312 299630 275324
rect 318794 275312 318800 275324
rect 299624 275284 318800 275312
rect 299624 275272 299630 275284
rect 318794 275272 318800 275284
rect 318852 275272 318858 275324
rect 297542 273912 297548 273964
rect 297600 273952 297606 273964
rect 335354 273952 335360 273964
rect 297600 273924 335360 273952
rect 297600 273912 297606 273924
rect 335354 273912 335360 273924
rect 335412 273912 335418 273964
rect 297634 273232 297640 273284
rect 297692 273272 297698 273284
rect 298738 273272 298744 273284
rect 297692 273244 298744 273272
rect 297692 273232 297698 273244
rect 298738 273232 298744 273244
rect 298796 273232 298802 273284
rect 479518 273164 479524 273216
rect 479576 273204 479582 273216
rect 579890 273204 579896 273216
rect 479576 273176 579896 273204
rect 479576 273164 479582 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 299658 271804 299664 271856
rect 299716 271844 299722 271856
rect 304994 271844 305000 271856
rect 299716 271816 305000 271844
rect 299716 271804 299722 271816
rect 304994 271804 305000 271816
rect 305052 271804 305058 271856
rect 13814 268404 13820 268456
rect 13872 268444 13878 268456
rect 485038 268444 485044 268456
rect 13872 268416 485044 268444
rect 13872 268404 13878 268416
rect 485038 268404 485044 268416
rect 485096 268404 485102 268456
rect 3418 268336 3424 268388
rect 3476 268376 3482 268388
rect 510982 268376 510988 268388
rect 3476 268348 510988 268376
rect 3476 268336 3482 268348
rect 510982 268336 510988 268348
rect 511040 268336 511046 268388
rect 301498 264188 301504 264240
rect 301556 264228 301562 264240
rect 350718 264228 350724 264240
rect 301556 264200 350724 264228
rect 301556 264188 301562 264200
rect 350718 264188 350724 264200
rect 350776 264188 350782 264240
rect 58986 262828 58992 262880
rect 59044 262868 59050 262880
rect 352374 262868 352380 262880
rect 59044 262840 352380 262868
rect 59044 262828 59050 262840
rect 352374 262828 352380 262840
rect 352432 262828 352438 262880
rect 58894 261468 58900 261520
rect 58952 261508 58958 261520
rect 352742 261508 352748 261520
rect 58952 261480 352748 261508
rect 58952 261468 58958 261480
rect 352742 261468 352748 261480
rect 352800 261468 352806 261520
rect 59262 260108 59268 260160
rect 59320 260148 59326 260160
rect 347866 260148 347872 260160
rect 59320 260120 347872 260148
rect 59320 260108 59326 260120
rect 347866 260108 347872 260120
rect 347924 260108 347930 260160
rect 356790 259360 356796 259412
rect 356848 259400 356854 259412
rect 579798 259400 579804 259412
rect 356848 259372 579804 259400
rect 356848 259360 356854 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 52454 250452 52460 250504
rect 52512 250492 52518 250504
rect 468570 250492 468576 250504
rect 52512 250464 468576 250492
rect 52512 250452 52518 250464
rect 468570 250452 468576 250464
rect 468628 250452 468634 250504
rect 359642 245556 359648 245608
rect 359700 245596 359706 245608
rect 580166 245596 580172 245608
rect 359700 245568 580172 245596
rect 359700 245556 359706 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3418 241408 3424 241460
rect 3476 241448 3482 241460
rect 510890 241448 510896 241460
rect 3476 241420 510896 241448
rect 3476 241408 3482 241420
rect 510890 241408 510896 241420
rect 510948 241408 510954 241460
rect 9674 239368 9680 239420
rect 9732 239408 9738 239420
rect 400858 239408 400864 239420
rect 9732 239380 400864 239408
rect 9732 239368 9738 239380
rect 400858 239368 400864 239380
rect 400916 239368 400922 239420
rect 59078 236648 59084 236700
rect 59136 236688 59142 236700
rect 352098 236688 352104 236700
rect 59136 236660 352104 236688
rect 59136 236648 59142 236660
rect 352098 236648 352104 236660
rect 352156 236648 352162 236700
rect 57054 233928 57060 233980
rect 57112 233968 57118 233980
rect 260282 233968 260288 233980
rect 57112 233940 260288 233968
rect 57112 233928 57118 233940
rect 260282 233928 260288 233940
rect 260340 233928 260346 233980
rect 14458 233860 14464 233912
rect 14516 233900 14522 233912
rect 490282 233900 490288 233912
rect 14516 233872 490288 233900
rect 14516 233860 14522 233872
rect 490282 233860 490288 233872
rect 490340 233860 490346 233912
rect 486418 233180 486424 233232
rect 486476 233220 486482 233232
rect 580166 233220 580172 233232
rect 486476 233192 580172 233220
rect 486476 233180 486482 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 59722 232500 59728 232552
rect 59780 232540 59786 232552
rect 311894 232540 311900 232552
rect 59780 232512 311900 232540
rect 59780 232500 59786 232512
rect 311894 232500 311900 232512
rect 311952 232500 311958 232552
rect 59630 229712 59636 229764
rect 59688 229752 59694 229764
rect 324406 229752 324412 229764
rect 59688 229724 324412 229752
rect 59688 229712 59694 229724
rect 324406 229712 324412 229724
rect 324464 229712 324470 229764
rect 325694 229712 325700 229764
rect 325752 229752 325758 229764
rect 349798 229752 349804 229764
rect 325752 229724 349804 229752
rect 325752 229712 325758 229724
rect 349798 229712 349804 229724
rect 349856 229712 349862 229764
rect 57422 228352 57428 228404
rect 57480 228392 57486 228404
rect 258718 228392 258724 228404
rect 57480 228364 258724 228392
rect 57480 228352 57486 228364
rect 258718 228352 258724 228364
rect 258776 228352 258782 228404
rect 59170 227060 59176 227112
rect 59228 227100 59234 227112
rect 283190 227100 283196 227112
rect 59228 227072 283196 227100
rect 59228 227060 59234 227072
rect 283190 227060 283196 227072
rect 283248 227060 283254 227112
rect 308858 227060 308864 227112
rect 308916 227100 308922 227112
rect 332594 227100 332600 227112
rect 308916 227072 332600 227100
rect 308916 227060 308922 227072
rect 332594 227060 332600 227072
rect 332652 227060 332658 227112
rect 57698 226992 57704 227044
rect 57756 227032 57762 227044
rect 293402 227032 293408 227044
rect 57756 227004 293408 227032
rect 57756 226992 57762 227004
rect 293402 226992 293408 227004
rect 293460 226992 293466 227044
rect 318978 226992 318984 227044
rect 319036 227032 319042 227044
rect 349706 227032 349712 227044
rect 319036 227004 349712 227032
rect 319036 226992 319042 227004
rect 349706 226992 349712 227004
rect 349764 226992 349770 227044
rect 302786 225768 302792 225820
rect 302844 225808 302850 225820
rect 381538 225808 381544 225820
rect 302844 225780 381544 225808
rect 302844 225768 302850 225780
rect 381538 225768 381544 225780
rect 381596 225768 381602 225820
rect 58802 225700 58808 225752
rect 58860 225740 58866 225752
rect 310606 225740 310612 225752
rect 58860 225712 310612 225740
rect 58860 225700 58866 225712
rect 310606 225700 310612 225712
rect 310664 225700 310670 225752
rect 42794 225632 42800 225684
rect 42852 225672 42858 225684
rect 512362 225672 512368 225684
rect 42852 225644 512368 225672
rect 42852 225632 42858 225644
rect 512362 225632 512368 225644
rect 512420 225632 512426 225684
rect 3510 225564 3516 225616
rect 3568 225604 3574 225616
rect 476942 225604 476948 225616
rect 3568 225576 476948 225604
rect 3568 225564 3574 225576
rect 476942 225564 476948 225576
rect 477000 225564 477006 225616
rect 3418 224272 3424 224324
rect 3476 224312 3482 224324
rect 436830 224312 436836 224324
rect 3476 224284 436836 224312
rect 3476 224272 3482 224284
rect 436830 224272 436836 224284
rect 436888 224272 436894 224324
rect 3694 224204 3700 224256
rect 3752 224244 3758 224256
rect 509878 224244 509884 224256
rect 3752 224216 509884 224244
rect 3752 224204 3758 224216
rect 509878 224204 509884 224216
rect 509936 224204 509942 224256
rect 305638 223524 305644 223576
rect 305696 223564 305702 223576
rect 307846 223564 307852 223576
rect 305696 223536 307852 223564
rect 305696 223524 305702 223536
rect 307846 223524 307852 223536
rect 307904 223524 307910 223576
rect 311158 223524 311164 223576
rect 311216 223564 311222 223576
rect 312906 223564 312912 223576
rect 311216 223536 312912 223564
rect 311216 223524 311222 223536
rect 312906 223524 312912 223536
rect 312964 223524 312970 223576
rect 326338 223524 326344 223576
rect 326396 223564 326402 223576
rect 333146 223564 333152 223576
rect 326396 223536 333152 223564
rect 326396 223524 326402 223536
rect 333146 223524 333152 223536
rect 333204 223524 333210 223576
rect 300118 223456 300124 223508
rect 300176 223496 300182 223508
rect 306834 223496 306840 223508
rect 300176 223468 306840 223496
rect 300176 223456 300182 223468
rect 306834 223456 306840 223468
rect 306892 223456 306898 223508
rect 335170 223252 335176 223304
rect 335228 223292 335234 223304
rect 341518 223292 341524 223304
rect 335228 223264 341524 223292
rect 335228 223252 335234 223264
rect 341518 223252 341524 223264
rect 341576 223252 341582 223304
rect 302234 223184 302240 223236
rect 302292 223224 302298 223236
rect 314930 223224 314936 223236
rect 302292 223196 314936 223224
rect 302292 223184 302298 223196
rect 314930 223184 314936 223196
rect 314988 223184 314994 223236
rect 337194 223184 337200 223236
rect 337252 223224 337258 223236
rect 349982 223224 349988 223236
rect 337252 223196 349988 223224
rect 337252 223184 337258 223196
rect 349982 223184 349988 223196
rect 350040 223184 350046 223236
rect 309226 223116 309232 223168
rect 309284 223156 309290 223168
rect 323026 223156 323032 223168
rect 309284 223128 323032 223156
rect 309284 223116 309290 223128
rect 323026 223116 323032 223128
rect 323084 223116 323090 223168
rect 329098 223116 329104 223168
rect 329156 223156 329162 223168
rect 354674 223156 354680 223168
rect 329156 223128 354680 223156
rect 329156 223116 329162 223128
rect 354674 223116 354680 223128
rect 354732 223116 354738 223168
rect 299750 223048 299756 223100
rect 299808 223088 299814 223100
rect 321002 223088 321008 223100
rect 299808 223060 321008 223088
rect 299808 223048 299814 223060
rect 321002 223048 321008 223060
rect 321060 223048 321066 223100
rect 328086 223048 328092 223100
rect 328144 223088 328150 223100
rect 353570 223088 353576 223100
rect 328144 223060 353576 223088
rect 328144 223048 328150 223060
rect 353570 223048 353576 223060
rect 353628 223048 353634 223100
rect 293862 222980 293868 223032
rect 293920 223020 293926 223032
rect 331122 223020 331128 223032
rect 293920 222992 331128 223020
rect 293920 222980 293926 222992
rect 331122 222980 331128 222992
rect 331180 222980 331186 223032
rect 334158 222980 334164 223032
rect 334216 223020 334222 223032
rect 354766 223020 354772 223032
rect 334216 222992 354772 223020
rect 334216 222980 334222 222992
rect 354766 222980 354772 222992
rect 354824 222980 354830 223032
rect 57790 222912 57796 222964
rect 57848 222952 57854 222964
rect 253566 222952 253572 222964
rect 57848 222924 253572 222952
rect 57848 222912 57854 222924
rect 253566 222912 253572 222924
rect 253624 222912 253630 222964
rect 293770 222912 293776 222964
rect 293828 222952 293834 222964
rect 311894 222952 311900 222964
rect 293828 222924 311900 222952
rect 293828 222912 293834 222924
rect 311894 222912 311900 222924
rect 311952 222912 311958 222964
rect 316954 222912 316960 222964
rect 317012 222952 317018 222964
rect 351362 222952 351368 222964
rect 317012 222924 351368 222952
rect 317012 222912 317018 222924
rect 351362 222912 351368 222924
rect 351420 222912 351426 222964
rect 57330 222844 57336 222896
rect 57388 222884 57394 222896
rect 254578 222884 254584 222896
rect 57388 222856 254584 222884
rect 57388 222844 57394 222856
rect 254578 222844 254584 222856
rect 254636 222844 254642 222896
rect 293678 222844 293684 222896
rect 293736 222884 293742 222896
rect 330110 222884 330116 222896
rect 293736 222856 330116 222884
rect 293736 222844 293742 222856
rect 330110 222844 330116 222856
rect 330168 222844 330174 222896
rect 332134 222844 332140 222896
rect 332192 222884 332198 222896
rect 353662 222884 353668 222896
rect 332192 222856 353668 222884
rect 332192 222844 332198 222856
rect 353662 222844 353668 222856
rect 353720 222844 353726 222896
rect 222838 222232 222844 222284
rect 222896 222272 222902 222284
rect 301498 222272 301504 222284
rect 222896 222244 301504 222272
rect 222896 222232 222902 222244
rect 301498 222232 301504 222244
rect 301556 222232 301562 222284
rect 224402 222164 224408 222216
rect 224460 222204 224466 222216
rect 339218 222204 339224 222216
rect 224460 222176 339224 222204
rect 224460 222164 224466 222176
rect 339218 222164 339224 222176
rect 339276 222164 339282 222216
rect 299474 222096 299480 222148
rect 299532 222136 299538 222148
rect 300762 222136 300768 222148
rect 299532 222108 300768 222136
rect 299532 222096 299538 222108
rect 300762 222096 300768 222108
rect 300820 222096 300826 222148
rect 298922 221552 298928 221604
rect 298980 221592 298986 221604
rect 313366 221592 313372 221604
rect 298980 221564 313372 221592
rect 298980 221552 298986 221564
rect 313366 221552 313372 221564
rect 313424 221552 313430 221604
rect 57238 221484 57244 221536
rect 57296 221524 57302 221536
rect 253382 221524 253388 221536
rect 57296 221496 253388 221524
rect 57296 221484 57302 221496
rect 253382 221484 253388 221496
rect 253440 221484 253446 221536
rect 297358 221484 297364 221536
rect 297416 221524 297422 221536
rect 337378 221524 337384 221536
rect 297416 221496 337384 221524
rect 297416 221484 297422 221496
rect 337378 221484 337384 221496
rect 337436 221484 337442 221536
rect 59814 221416 59820 221468
rect 59872 221456 59878 221468
rect 352282 221456 352288 221468
rect 59872 221428 352288 221456
rect 59872 221416 59878 221428
rect 352282 221416 352288 221428
rect 352340 221416 352346 221468
rect 226058 220804 226064 220856
rect 226116 220844 226122 220856
rect 300762 220844 300768 220856
rect 226116 220816 300768 220844
rect 226116 220804 226122 220816
rect 300762 220804 300768 220816
rect 300820 220844 300826 220856
rect 578878 220844 578884 220856
rect 300820 220816 578884 220844
rect 300820 220804 300826 220816
rect 578878 220804 578884 220816
rect 578936 220804 578942 220856
rect 299014 220260 299020 220312
rect 299072 220300 299078 220312
rect 306374 220300 306380 220312
rect 299072 220272 306380 220300
rect 299072 220260 299078 220272
rect 306374 220260 306380 220272
rect 306432 220260 306438 220312
rect 57146 220192 57152 220244
rect 57204 220232 57210 220244
rect 291930 220232 291936 220244
rect 57204 220204 291936 220232
rect 57204 220192 57210 220204
rect 291930 220192 291936 220204
rect 291988 220192 291994 220244
rect 298830 220192 298836 220244
rect 298888 220232 298894 220244
rect 328454 220232 328460 220244
rect 298888 220204 328460 220232
rect 298888 220192 298894 220204
rect 328454 220192 328460 220204
rect 328512 220192 328518 220244
rect 60550 220124 60556 220176
rect 60608 220164 60614 220176
rect 294598 220164 294604 220176
rect 60608 220136 294604 220164
rect 60608 220124 60614 220136
rect 294598 220124 294604 220136
rect 294656 220124 294662 220176
rect 297266 220124 297272 220176
rect 297324 220164 297330 220176
rect 336918 220164 336924 220176
rect 297324 220136 336924 220164
rect 297324 220124 297330 220136
rect 336918 220124 336924 220136
rect 336976 220124 336982 220176
rect 3602 220056 3608 220108
rect 3660 220096 3666 220108
rect 510798 220096 510804 220108
rect 3660 220068 510804 220096
rect 3660 220056 3666 220068
rect 510798 220056 510804 220068
rect 510856 220056 510862 220108
rect 351270 219376 351276 219428
rect 351328 219416 351334 219428
rect 579890 219416 579896 219428
rect 351328 219388 579896 219416
rect 351328 219376 351334 219388
rect 579890 219376 579896 219388
rect 579948 219376 579954 219428
rect 57882 218764 57888 218816
rect 57940 218804 57946 218816
rect 253198 218804 253204 218816
rect 57940 218776 253204 218804
rect 57940 218764 57946 218776
rect 253198 218764 253204 218776
rect 253256 218764 253262 218816
rect 57606 218696 57612 218748
rect 57664 218736 57670 218748
rect 293218 218736 293224 218748
rect 57664 218708 293224 218736
rect 57664 218696 57670 218708
rect 293218 218696 293224 218708
rect 293276 218696 293282 218748
rect 222930 216656 222936 216708
rect 222988 216696 222994 216708
rect 296806 216696 296812 216708
rect 222988 216668 296812 216696
rect 222988 216656 222994 216668
rect 296806 216656 296812 216668
rect 296864 216656 296870 216708
rect 247678 215296 247684 215348
rect 247736 215336 247742 215348
rect 297726 215336 297732 215348
rect 247736 215308 297732 215336
rect 247736 215296 247742 215308
rect 297726 215296 297732 215308
rect 297784 215296 297790 215348
rect 57238 214548 57244 214600
rect 57296 214588 57302 214600
rect 57514 214588 57520 214600
rect 57296 214560 57520 214588
rect 57296 214548 57302 214560
rect 57514 214548 57520 214560
rect 57572 214548 57578 214600
rect 246298 213936 246304 213988
rect 246356 213976 246362 213988
rect 297726 213976 297732 213988
rect 246356 213948 297732 213976
rect 246356 213936 246362 213948
rect 297726 213936 297732 213948
rect 297784 213936 297790 213988
rect 222286 212984 222292 213036
rect 222344 213024 222350 213036
rect 226058 213024 226064 213036
rect 222344 212996 226064 213024
rect 222344 212984 222350 212996
rect 226058 212984 226064 212996
rect 226116 212984 226122 213036
rect 243538 212508 243544 212560
rect 243596 212548 243602 212560
rect 297726 212548 297732 212560
rect 243596 212520 297732 212548
rect 243596 212508 243602 212520
rect 297726 212508 297732 212520
rect 297784 212508 297790 212560
rect 242158 211148 242164 211200
rect 242216 211188 242222 211200
rect 297726 211188 297732 211200
rect 242216 211160 297732 211188
rect 242216 211148 242222 211160
rect 297726 211148 297732 211160
rect 297784 211148 297790 211200
rect 239398 209788 239404 209840
rect 239456 209828 239462 209840
rect 297726 209828 297732 209840
rect 239456 209800 297732 209828
rect 239456 209788 239462 209800
rect 297726 209788 297732 209800
rect 297784 209788 297790 209840
rect 238018 208360 238024 208412
rect 238076 208400 238082 208412
rect 297726 208400 297732 208412
rect 238076 208372 297732 208400
rect 238076 208360 238082 208372
rect 297726 208360 297732 208372
rect 297784 208360 297790 208412
rect 232498 207000 232504 207052
rect 232556 207040 232562 207052
rect 297726 207040 297732 207052
rect 232556 207012 297732 207040
rect 232556 207000 232562 207012
rect 297726 207000 297732 207012
rect 297784 207000 297790 207052
rect 418798 206932 418804 206984
rect 418856 206972 418862 206984
rect 580166 206972 580172 206984
rect 418856 206944 580172 206972
rect 418856 206932 418862 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 229738 205640 229744 205692
rect 229796 205680 229802 205692
rect 297726 205680 297732 205692
rect 229796 205652 297732 205680
rect 229796 205640 229802 205652
rect 297726 205640 297732 205652
rect 297784 205640 297790 205692
rect 223206 205572 223212 205624
rect 223264 205612 223270 205624
rect 229830 205612 229836 205624
rect 223264 205584 229836 205612
rect 223264 205572 223270 205584
rect 229830 205572 229836 205584
rect 229888 205572 229894 205624
rect 287698 201492 287704 201544
rect 287756 201532 287762 201544
rect 296806 201532 296812 201544
rect 287756 201504 296812 201532
rect 287756 201492 287762 201504
rect 296806 201492 296812 201504
rect 296864 201492 296870 201544
rect 51718 201424 51724 201476
rect 51776 201464 51782 201476
rect 57330 201464 57336 201476
rect 51776 201436 57336 201464
rect 51776 201424 51782 201436
rect 57330 201424 57336 201436
rect 57388 201424 57394 201476
rect 228358 200132 228364 200184
rect 228416 200172 228422 200184
rect 297726 200172 297732 200184
rect 228416 200144 297732 200172
rect 228416 200132 228422 200144
rect 297726 200132 297732 200144
rect 297784 200132 297790 200184
rect 225598 198704 225604 198756
rect 225656 198744 225662 198756
rect 297726 198744 297732 198756
rect 225656 198716 297732 198744
rect 225656 198704 225662 198716
rect 297726 198704 297732 198716
rect 297784 198704 297790 198756
rect 224310 197344 224316 197396
rect 224368 197384 224374 197396
rect 297726 197384 297732 197396
rect 224368 197356 297732 197384
rect 224368 197344 224374 197356
rect 297726 197344 297732 197356
rect 297784 197344 297790 197396
rect 50982 197276 50988 197328
rect 51040 197316 51046 197328
rect 57330 197316 57336 197328
rect 51040 197288 57336 197316
rect 51040 197276 51046 197288
rect 57330 197276 57336 197288
rect 57388 197276 57394 197328
rect 224218 195984 224224 196036
rect 224276 196024 224282 196036
rect 297726 196024 297732 196036
rect 224276 195996 297732 196024
rect 224276 195984 224282 195996
rect 297726 195984 297732 195996
rect 297784 195984 297790 196036
rect 223482 194556 223488 194608
rect 223540 194596 223546 194608
rect 233970 194596 233976 194608
rect 223540 194568 233976 194596
rect 223540 194556 223546 194568
rect 233970 194556 233976 194568
rect 234028 194556 234034 194608
rect 250438 194556 250444 194608
rect 250496 194596 250502 194608
rect 297726 194596 297732 194608
rect 250496 194568 297732 194596
rect 250496 194556 250502 194568
rect 297726 194556 297732 194568
rect 297784 194556 297790 194608
rect 235258 193196 235264 193248
rect 235316 193236 235322 193248
rect 297726 193236 297732 193248
rect 235316 193208 297732 193236
rect 235316 193196 235322 193208
rect 297726 193196 297732 193208
rect 297784 193196 297790 193248
rect 229830 193128 229836 193180
rect 229888 193168 229894 193180
rect 297542 193168 297548 193180
rect 229888 193140 297548 193168
rect 229888 193128 229894 193140
rect 297542 193128 297548 193140
rect 297600 193128 297606 193180
rect 552658 193128 552664 193180
rect 552716 193168 552722 193180
rect 580166 193168 580172 193180
rect 552716 193140 580172 193168
rect 552716 193128 552722 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 50890 192448 50896 192500
rect 50948 192488 50954 192500
rect 57238 192488 57244 192500
rect 50948 192460 57244 192488
rect 50948 192448 50954 192460
rect 57238 192448 57244 192460
rect 57296 192448 57302 192500
rect 223482 191836 223488 191888
rect 223540 191876 223546 191888
rect 229922 191876 229928 191888
rect 223540 191848 229928 191876
rect 223540 191836 223546 191848
rect 229922 191836 229928 191848
rect 229980 191836 229986 191888
rect 233878 190476 233884 190528
rect 233936 190516 233942 190528
rect 297726 190516 297732 190528
rect 233936 190488 297732 190516
rect 233936 190476 233942 190488
rect 297726 190476 297732 190488
rect 297784 190476 297790 190528
rect 222838 190408 222844 190460
rect 222896 190448 222902 190460
rect 297542 190448 297548 190460
rect 222896 190420 297548 190448
rect 222896 190408 222902 190420
rect 297542 190408 297548 190420
rect 297600 190408 297606 190460
rect 222838 189048 222844 189100
rect 222896 189088 222902 189100
rect 224954 189088 224960 189100
rect 222896 189060 224960 189088
rect 222896 189048 222902 189060
rect 224954 189048 224960 189060
rect 225012 189048 225018 189100
rect 50430 188980 50436 189032
rect 50488 189020 50494 189032
rect 57330 189020 57336 189032
rect 50488 188992 57336 189020
rect 50488 188980 50494 188992
rect 57330 188980 57336 188992
rect 57388 188980 57394 189032
rect 223022 188980 223028 189032
rect 223080 189020 223086 189032
rect 297726 189020 297732 189032
rect 223080 188992 297732 189020
rect 223080 188980 223086 188992
rect 297726 188980 297732 188992
rect 297784 188980 297790 189032
rect 222838 186328 222844 186380
rect 222896 186368 222902 186380
rect 228450 186368 228456 186380
rect 222896 186340 228456 186368
rect 222896 186328 222902 186340
rect 228450 186328 228456 186340
rect 228508 186328 228514 186380
rect 222930 186260 222936 186312
rect 222988 186300 222994 186312
rect 297726 186300 297732 186312
rect 222988 186272 297732 186300
rect 222988 186260 222994 186272
rect 297726 186260 297732 186272
rect 297784 186260 297790 186312
rect 51074 184832 51080 184884
rect 51132 184872 51138 184884
rect 56686 184872 56692 184884
rect 51132 184844 56692 184872
rect 51132 184832 51138 184844
rect 56686 184832 56692 184844
rect 56744 184832 56750 184884
rect 233970 184832 233976 184884
rect 234028 184872 234034 184884
rect 297726 184872 297732 184884
rect 234028 184844 297732 184872
rect 234028 184832 234034 184844
rect 297726 184832 297732 184844
rect 297784 184832 297790 184884
rect 222286 183744 222292 183796
rect 222344 183784 222350 183796
rect 225782 183784 225788 183796
rect 222344 183756 225788 183784
rect 222344 183744 222350 183756
rect 225782 183744 225788 183756
rect 225840 183744 225846 183796
rect 229922 183472 229928 183524
rect 229980 183512 229986 183524
rect 297726 183512 297732 183524
rect 229980 183484 297732 183512
rect 229980 183472 229986 183484
rect 297726 183472 297732 183484
rect 297784 183472 297790 183524
rect 224954 182112 224960 182164
rect 225012 182152 225018 182164
rect 297726 182152 297732 182164
rect 225012 182124 297732 182152
rect 225012 182112 225018 182124
rect 297726 182112 297732 182124
rect 297784 182112 297790 182164
rect 51166 180752 51172 180804
rect 51224 180792 51230 180804
rect 56686 180792 56692 180804
rect 51224 180764 56692 180792
rect 51224 180752 51230 180764
rect 56686 180752 56692 180764
rect 56744 180752 56750 180804
rect 228450 180752 228456 180804
rect 228508 180792 228514 180804
rect 297726 180792 297732 180804
rect 228508 180764 297732 180792
rect 228508 180752 228514 180764
rect 297726 180752 297732 180764
rect 297784 180752 297790 180804
rect 225782 179324 225788 179376
rect 225840 179364 225846 179376
rect 297726 179364 297732 179376
rect 225840 179336 297732 179364
rect 225840 179324 225846 179336
rect 297726 179324 297732 179336
rect 297784 179324 297790 179376
rect 223482 177964 223488 178016
rect 223540 178004 223546 178016
rect 297726 178004 297732 178016
rect 223540 177976 297732 178004
rect 223540 177964 223546 177976
rect 297726 177964 297732 177976
rect 297784 177964 297790 178016
rect 477862 177352 477868 177404
rect 477920 177392 477926 177404
rect 516134 177392 516140 177404
rect 477920 177364 516140 177392
rect 477920 177352 477926 177364
rect 516134 177352 516140 177364
rect 516192 177352 516198 177404
rect 358446 177284 358452 177336
rect 358504 177324 358510 177336
rect 426434 177324 426440 177336
rect 358504 177296 426440 177324
rect 358504 177284 358510 177296
rect 426434 177284 426440 177296
rect 426492 177284 426498 177336
rect 478506 177284 478512 177336
rect 478564 177324 478570 177336
rect 520274 177324 520280 177336
rect 478564 177296 520280 177324
rect 478564 177284 478570 177296
rect 520274 177284 520280 177296
rect 520332 177284 520338 177336
rect 50338 176604 50344 176656
rect 50396 176644 50402 176656
rect 57330 176644 57336 176656
rect 50396 176616 57336 176644
rect 50396 176604 50402 176616
rect 57330 176604 57336 176616
rect 57388 176604 57394 176656
rect 222654 176604 222660 176656
rect 222712 176644 222718 176656
rect 297726 176644 297732 176656
rect 222712 176616 297732 176644
rect 222712 176604 222718 176616
rect 297726 176604 297732 176616
rect 297784 176604 297790 176656
rect 222654 175176 222660 175228
rect 222712 175216 222718 175228
rect 297726 175216 297732 175228
rect 222712 175188 297732 175216
rect 222712 175176 222718 175188
rect 297726 175176 297732 175188
rect 297784 175176 297790 175228
rect 48866 173340 48872 173392
rect 48924 173380 48930 173392
rect 57238 173380 57244 173392
rect 48924 173352 57244 173380
rect 48924 173340 48930 173352
rect 57238 173340 57244 173352
rect 57296 173340 57302 173392
rect 222378 173136 222384 173188
rect 222436 173176 222442 173188
rect 297726 173176 297732 173188
rect 222436 173148 297732 173176
rect 222436 173136 222442 173148
rect 297726 173136 297732 173148
rect 297784 173136 297790 173188
rect 222470 171096 222476 171148
rect 222528 171136 222534 171148
rect 297726 171136 297732 171148
rect 222528 171108 297732 171136
rect 222528 171096 222534 171108
rect 297726 171096 297732 171108
rect 297784 171096 297790 171148
rect 222930 169736 222936 169788
rect 222988 169776 222994 169788
rect 297726 169776 297732 169788
rect 222988 169748 297732 169776
rect 222988 169736 222994 169748
rect 297726 169736 297732 169748
rect 297784 169736 297790 169788
rect 49510 169668 49516 169720
rect 49568 169708 49574 169720
rect 57330 169708 57336 169720
rect 49568 169680 57336 169708
rect 49568 169668 49574 169680
rect 57330 169668 57336 169680
rect 57388 169668 57394 169720
rect 223482 167016 223488 167068
rect 223540 167056 223546 167068
rect 297726 167056 297732 167068
rect 223540 167028 297732 167056
rect 223540 167016 223546 167028
rect 297726 167016 297732 167028
rect 297784 167016 297790 167068
rect 409138 166948 409144 167000
rect 409196 166988 409202 167000
rect 580166 166988 580172 167000
rect 409196 166960 580172 166988
rect 409196 166948 409202 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 223022 165588 223028 165640
rect 223080 165628 223086 165640
rect 296806 165628 296812 165640
rect 223080 165600 296812 165628
rect 223080 165588 223086 165600
rect 296806 165588 296812 165600
rect 296864 165588 296870 165640
rect 222930 164228 222936 164280
rect 222988 164268 222994 164280
rect 297726 164268 297732 164280
rect 222988 164240 297732 164268
rect 222988 164228 222994 164240
rect 297726 164228 297732 164240
rect 297784 164228 297790 164280
rect 223482 162868 223488 162920
rect 223540 162908 223546 162920
rect 297726 162908 297732 162920
rect 223540 162880 297732 162908
rect 223540 162868 223546 162880
rect 297726 162868 297732 162880
rect 297784 162868 297790 162920
rect 229094 161440 229100 161492
rect 229152 161480 229158 161492
rect 297726 161480 297732 161492
rect 229152 161452 297732 161480
rect 229152 161440 229158 161452
rect 297726 161440 297732 161452
rect 297784 161440 297790 161492
rect 54570 161372 54576 161424
rect 54628 161412 54634 161424
rect 57054 161412 57060 161424
rect 54628 161384 57060 161412
rect 54628 161372 54634 161384
rect 57054 161372 57060 161384
rect 57112 161372 57118 161424
rect 231118 160080 231124 160132
rect 231176 160120 231182 160132
rect 297726 160120 297732 160132
rect 231176 160092 297732 160120
rect 231176 160080 231182 160092
rect 297726 160080 297732 160092
rect 297784 160080 297790 160132
rect 228450 158720 228456 158772
rect 228508 158760 228514 158772
rect 297726 158760 297732 158772
rect 228508 158732 297732 158760
rect 228508 158720 228514 158732
rect 297726 158720 297732 158732
rect 297784 158720 297790 158772
rect 225690 157360 225696 157412
rect 225748 157400 225754 157412
rect 296806 157400 296812 157412
rect 225748 157372 296812 157400
rect 225748 157360 225754 157372
rect 296806 157360 296812 157372
rect 296864 157360 296870 157412
rect 53098 157292 53104 157344
rect 53156 157332 53162 157344
rect 57054 157332 57060 157344
rect 53156 157304 57060 157332
rect 53156 157292 53162 157304
rect 57054 157292 57060 157304
rect 57112 157292 57118 157344
rect 222562 157088 222568 157140
rect 222620 157128 222626 157140
rect 229094 157128 229100 157140
rect 222620 157100 229100 157128
rect 222620 157088 222626 157100
rect 229094 157088 229100 157100
rect 229152 157088 229158 157140
rect 229830 155932 229836 155984
rect 229888 155972 229894 155984
rect 297726 155972 297732 155984
rect 229888 155944 297732 155972
rect 229888 155932 229894 155944
rect 297726 155932 297732 155944
rect 297784 155932 297790 155984
rect 222930 154572 222936 154624
rect 222988 154612 222994 154624
rect 297726 154612 297732 154624
rect 222988 154584 297732 154612
rect 222988 154572 222994 154584
rect 297726 154572 297732 154584
rect 297784 154572 297790 154624
rect 222838 153212 222844 153264
rect 222896 153252 222902 153264
rect 297726 153252 297732 153264
rect 222896 153224 297732 153252
rect 222896 153212 222902 153224
rect 297726 153212 297732 153224
rect 297784 153212 297790 153264
rect 54478 153144 54484 153196
rect 54536 153184 54542 153196
rect 57330 153184 57336 153196
rect 54536 153156 57336 153184
rect 54536 153144 54542 153156
rect 57330 153144 57336 153156
rect 57388 153144 57394 153196
rect 536098 153144 536104 153196
rect 536156 153184 536162 153196
rect 579798 153184 579804 153196
rect 536156 153156 579804 153184
rect 536156 153144 536162 153156
rect 579798 153144 579804 153156
rect 579856 153144 579862 153196
rect 236638 151784 236644 151836
rect 236696 151824 236702 151836
rect 297726 151824 297732 151836
rect 236696 151796 297732 151824
rect 236696 151784 236702 151796
rect 297726 151784 297732 151796
rect 297784 151784 297790 151836
rect 223482 150424 223488 150476
rect 223540 150464 223546 150476
rect 231118 150464 231124 150476
rect 223540 150436 231124 150464
rect 223540 150424 223546 150436
rect 231118 150424 231124 150436
rect 231176 150424 231182 150476
rect 235350 149064 235356 149116
rect 235408 149104 235414 149116
rect 297726 149104 297732 149116
rect 235408 149076 297732 149104
rect 235408 149064 235414 149076
rect 297726 149064 297732 149076
rect 297784 149064 297790 149116
rect 50798 148996 50804 149048
rect 50856 149036 50862 149048
rect 57330 149036 57336 149048
rect 50856 149008 57336 149036
rect 50856 148996 50862 149008
rect 57330 148996 57336 149008
rect 57388 148996 57394 149048
rect 233970 147636 233976 147688
rect 234028 147676 234034 147688
rect 296806 147676 296812 147688
rect 234028 147648 296812 147676
rect 234028 147636 234034 147648
rect 296806 147636 296812 147648
rect 296864 147636 296870 147688
rect 223482 147228 223488 147280
rect 223540 147268 223546 147280
rect 228450 147268 228456 147280
rect 223540 147240 228456 147268
rect 223540 147228 223546 147240
rect 228450 147228 228456 147240
rect 228508 147228 228514 147280
rect 231118 146276 231124 146328
rect 231176 146316 231182 146328
rect 297726 146316 297732 146328
rect 231176 146288 297732 146316
rect 231176 146276 231182 146288
rect 297726 146276 297732 146288
rect 297784 146276 297790 146328
rect 228450 144916 228456 144968
rect 228508 144956 228514 144968
rect 297726 144956 297732 144968
rect 228508 144928 297732 144956
rect 228508 144916 228514 144928
rect 297726 144916 297732 144928
rect 297784 144916 297790 144968
rect 50706 144508 50712 144560
rect 50764 144548 50770 144560
rect 57330 144548 57336 144560
rect 50764 144520 57336 144548
rect 50764 144508 50770 144520
rect 57330 144508 57336 144520
rect 57388 144508 57394 144560
rect 222470 144304 222476 144356
rect 222528 144344 222534 144356
rect 225690 144344 225696 144356
rect 222528 144316 225696 144344
rect 222528 144304 222534 144316
rect 225690 144304 225696 144316
rect 225748 144304 225754 144356
rect 232590 143556 232596 143608
rect 232648 143596 232654 143608
rect 297726 143596 297732 143608
rect 232648 143568 297732 143596
rect 232648 143556 232654 143568
rect 297726 143556 297732 143568
rect 297784 143556 297790 143608
rect 251818 142128 251824 142180
rect 251876 142168 251882 142180
rect 297542 142168 297548 142180
rect 251876 142140 297548 142168
rect 251876 142128 251882 142140
rect 297542 142128 297548 142140
rect 297600 142128 297606 142180
rect 257338 142060 257344 142112
rect 257396 142100 257402 142112
rect 297726 142100 297732 142112
rect 257396 142072 297732 142100
rect 257396 142060 257402 142072
rect 297726 142060 297732 142072
rect 297784 142060 297790 142112
rect 223482 141448 223488 141500
rect 223540 141488 223546 141500
rect 229830 141488 229836 141500
rect 223540 141460 229836 141488
rect 223540 141448 223546 141460
rect 229830 141448 229836 141460
rect 229888 141448 229894 141500
rect 51258 140700 51264 140752
rect 51316 140740 51322 140752
rect 57422 140740 57428 140752
rect 51316 140712 57428 140740
rect 51316 140700 51322 140712
rect 57422 140700 57428 140712
rect 57480 140700 57486 140752
rect 273990 140700 273996 140752
rect 274048 140740 274054 140752
rect 297726 140740 297732 140752
rect 274048 140712 297732 140740
rect 274048 140700 274054 140712
rect 297726 140700 297732 140712
rect 297784 140700 297790 140752
rect 271230 139340 271236 139392
rect 271288 139380 271294 139392
rect 297726 139380 297732 139392
rect 271288 139352 297732 139380
rect 271288 139340 271294 139352
rect 297726 139340 297732 139352
rect 297784 139340 297790 139392
rect 353938 139340 353944 139392
rect 353996 139380 354002 139392
rect 580166 139380 580172 139392
rect 353996 139352 580172 139380
rect 353996 139340 354002 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 278038 137912 278044 137964
rect 278096 137952 278102 137964
rect 297726 137952 297732 137964
rect 278096 137924 297732 137952
rect 278096 137912 278102 137924
rect 297726 137912 297732 137924
rect 297784 137912 297790 137964
rect 3142 137708 3148 137760
rect 3200 137748 3206 137760
rect 8938 137748 8944 137760
rect 3200 137720 8944 137748
rect 3200 137708 3206 137720
rect 8938 137708 8944 137720
rect 8996 137708 9002 137760
rect 222470 137232 222476 137284
rect 222528 137272 222534 137284
rect 236638 137272 236644 137284
rect 222528 137244 236644 137272
rect 222528 137232 222534 137244
rect 236638 137232 236644 137244
rect 236696 137232 236702 137284
rect 269850 136552 269856 136604
rect 269908 136592 269914 136604
rect 296806 136592 296812 136604
rect 269908 136564 296812 136592
rect 269908 136552 269914 136564
rect 296806 136552 296812 136564
rect 296864 136552 296870 136604
rect 275370 135192 275376 135244
rect 275428 135232 275434 135244
rect 297726 135232 297732 135244
rect 275428 135204 297732 135232
rect 275428 135192 275434 135204
rect 297726 135192 297732 135204
rect 297784 135192 297790 135244
rect 223114 133152 223120 133204
rect 223172 133192 223178 133204
rect 235350 133192 235356 133204
rect 223172 133164 235356 133192
rect 223172 133152 223178 133164
rect 235350 133152 235356 133164
rect 235408 133152 235414 133204
rect 274082 132404 274088 132456
rect 274140 132444 274146 132456
rect 297726 132444 297732 132456
rect 274140 132416 297732 132444
rect 274140 132404 274146 132416
rect 297726 132404 297732 132416
rect 297784 132404 297790 132456
rect 271322 131044 271328 131096
rect 271380 131084 271386 131096
rect 297726 131084 297732 131096
rect 271380 131056 297732 131084
rect 271380 131044 271386 131056
rect 297726 131044 297732 131056
rect 297784 131044 297790 131096
rect 223482 130364 223488 130416
rect 223540 130404 223546 130416
rect 233970 130404 233976 130416
rect 223540 130376 233976 130404
rect 223540 130364 223546 130376
rect 233970 130364 233976 130376
rect 234028 130364 234034 130416
rect 275462 129684 275468 129736
rect 275520 129724 275526 129736
rect 297726 129724 297732 129736
rect 275520 129696 297732 129724
rect 275520 129684 275526 129696
rect 297726 129684 297732 129696
rect 297784 129684 297790 129736
rect 222470 128256 222476 128308
rect 222528 128296 222534 128308
rect 231118 128296 231124 128308
rect 222528 128268 231124 128296
rect 222528 128256 222534 128268
rect 231118 128256 231124 128268
rect 231176 128256 231182 128308
rect 257430 128256 257436 128308
rect 257488 128296 257494 128308
rect 297726 128296 297732 128308
rect 257488 128268 297732 128296
rect 257488 128256 257494 128268
rect 297726 128256 297732 128268
rect 297784 128256 297790 128308
rect 261570 126896 261576 126948
rect 261628 126936 261634 126948
rect 297726 126936 297732 126948
rect 261628 126908 297732 126936
rect 261628 126896 261634 126908
rect 297726 126896 297732 126908
rect 297784 126896 297790 126948
rect 372890 126896 372896 126948
rect 372948 126936 372954 126948
rect 580166 126936 580172 126948
rect 372948 126908 580172 126936
rect 372948 126896 372954 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 279418 125536 279424 125588
rect 279476 125576 279482 125588
rect 297726 125576 297732 125588
rect 279476 125548 297732 125576
rect 279476 125536 279482 125548
rect 297726 125536 297732 125548
rect 297784 125536 297790 125588
rect 223206 124584 223212 124636
rect 223264 124624 223270 124636
rect 228450 124624 228456 124636
rect 223264 124596 228456 124624
rect 223264 124584 223270 124596
rect 228450 124584 228456 124596
rect 228508 124584 228514 124636
rect 268470 124108 268476 124160
rect 268528 124148 268534 124160
rect 297726 124148 297732 124160
rect 268528 124120 297732 124148
rect 268528 124108 268534 124120
rect 297726 124108 297732 124120
rect 297784 124108 297790 124160
rect 265710 122748 265716 122800
rect 265768 122788 265774 122800
rect 297726 122788 297732 122800
rect 265768 122760 297732 122788
rect 265768 122748 265774 122760
rect 297726 122748 297732 122760
rect 297784 122748 297790 122800
rect 264330 121388 264336 121440
rect 264388 121428 264394 121440
rect 297726 121428 297732 121440
rect 264388 121400 297732 121428
rect 264388 121388 264394 121400
rect 297726 121388 297732 121400
rect 297784 121388 297790 121440
rect 289078 120028 289084 120080
rect 289136 120068 289142 120080
rect 297726 120068 297732 120080
rect 289136 120040 297732 120068
rect 289136 120028 289142 120040
rect 297726 120028 297732 120040
rect 297784 120028 297790 120080
rect 223482 118600 223488 118652
rect 223540 118640 223546 118652
rect 232590 118640 232596 118652
rect 223540 118612 232596 118640
rect 223540 118600 223546 118612
rect 232590 118600 232596 118612
rect 232648 118600 232654 118652
rect 269942 118600 269948 118652
rect 270000 118640 270006 118652
rect 296806 118640 296812 118652
rect 270000 118612 296812 118640
rect 270000 118600 270006 118612
rect 296806 118600 296812 118612
rect 296864 118600 296870 118652
rect 284938 117240 284944 117292
rect 284996 117280 285002 117292
rect 297726 117280 297732 117292
rect 284996 117252 297732 117280
rect 284996 117240 285002 117252
rect 297726 117240 297732 117252
rect 297784 117240 297790 117292
rect 342898 117240 342904 117292
rect 342956 117280 342962 117292
rect 475562 117280 475568 117292
rect 342956 117252 475568 117280
rect 342956 117240 342962 117252
rect 475562 117240 475568 117252
rect 475620 117240 475626 117292
rect 223482 115880 223488 115932
rect 223540 115920 223546 115932
rect 251818 115920 251824 115932
rect 223540 115892 251824 115920
rect 223540 115880 223546 115892
rect 251818 115880 251824 115892
rect 251876 115880 251882 115932
rect 278222 114452 278228 114504
rect 278280 114492 278286 114504
rect 297726 114492 297732 114504
rect 278280 114464 297732 114492
rect 278280 114452 278286 114464
rect 297726 114452 297732 114464
rect 297784 114452 297790 114504
rect 257522 113092 257528 113144
rect 257580 113132 257586 113144
rect 297726 113132 297732 113144
rect 257580 113104 297732 113132
rect 257580 113092 257586 113104
rect 297726 113092 297732 113104
rect 297784 113092 297790 113144
rect 571978 113092 571984 113144
rect 572036 113132 572042 113144
rect 580166 113132 580172 113144
rect 572036 113104 580172 113132
rect 572036 113092 572042 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 222194 112956 222200 113008
rect 222252 112996 222258 113008
rect 224402 112996 224408 113008
rect 222252 112968 224408 112996
rect 222252 112956 222258 112968
rect 224402 112956 224408 112968
rect 224460 112956 224466 113008
rect 223482 110372 223488 110424
rect 223540 110412 223546 110424
rect 247678 110412 247684 110424
rect 223540 110384 247684 110412
rect 223540 110372 223546 110384
rect 247678 110372 247684 110384
rect 247736 110372 247742 110424
rect 342898 108944 342904 108996
rect 342956 108984 342962 108996
rect 481082 108984 481088 108996
rect 342956 108956 481088 108984
rect 342956 108944 342962 108956
rect 481082 108944 481088 108956
rect 481140 108944 481146 108996
rect 222654 107584 222660 107636
rect 222712 107624 222718 107636
rect 246298 107624 246304 107636
rect 222712 107596 246304 107624
rect 222712 107584 222718 107596
rect 246298 107584 246304 107596
rect 246356 107584 246362 107636
rect 342898 106224 342904 106276
rect 342956 106264 342962 106276
rect 505094 106264 505100 106276
rect 342956 106236 505100 106264
rect 342956 106224 342962 106236
rect 505094 106224 505100 106236
rect 505152 106224 505158 106276
rect 222838 104796 222844 104848
rect 222896 104836 222902 104848
rect 243538 104836 243544 104848
rect 222896 104808 243544 104836
rect 222896 104796 222902 104808
rect 243538 104796 243544 104808
rect 243596 104796 243602 104848
rect 223482 102076 223488 102128
rect 223540 102116 223546 102128
rect 242158 102116 242164 102128
rect 223540 102088 242164 102116
rect 223540 102076 223546 102088
rect 242158 102076 242164 102088
rect 242216 102076 242222 102128
rect 223022 99288 223028 99340
rect 223080 99328 223086 99340
rect 239398 99328 239404 99340
rect 223080 99300 239404 99328
rect 223080 99288 223086 99300
rect 239398 99288 239404 99300
rect 239456 99288 239462 99340
rect 223114 96568 223120 96620
rect 223172 96608 223178 96620
rect 238018 96608 238024 96620
rect 223172 96580 238024 96608
rect 223172 96568 223178 96580
rect 238018 96568 238024 96580
rect 238076 96568 238082 96620
rect 223482 93780 223488 93832
rect 223540 93820 223546 93832
rect 232498 93820 232504 93832
rect 223540 93792 232504 93820
rect 223540 93780 223546 93792
rect 232498 93780 232504 93792
rect 232556 93780 232562 93832
rect 223390 91740 223396 91792
rect 223448 91780 223454 91792
rect 295978 91780 295984 91792
rect 223448 91752 295984 91780
rect 223448 91740 223454 91752
rect 295978 91740 295984 91752
rect 296036 91740 296042 91792
rect 223482 90312 223488 90364
rect 223540 90352 223546 90364
rect 229738 90352 229744 90364
rect 223540 90324 229744 90352
rect 223540 90312 223546 90324
rect 229738 90312 229744 90324
rect 229796 90312 229802 90364
rect 264238 90312 264244 90364
rect 264296 90352 264302 90364
rect 296806 90352 296812 90364
rect 264296 90324 296812 90352
rect 264296 90312 264302 90324
rect 296806 90312 296812 90324
rect 296864 90312 296870 90364
rect 358538 89020 358544 89072
rect 358596 89060 358602 89072
rect 408494 89060 408500 89072
rect 358596 89032 408500 89060
rect 358596 89020 358602 89032
rect 408494 89020 408500 89032
rect 408552 89020 408558 89072
rect 260190 88952 260196 89004
rect 260248 88992 260254 89004
rect 297358 88992 297364 89004
rect 260248 88964 297364 88992
rect 260248 88952 260254 88964
rect 297358 88952 297364 88964
rect 297416 88952 297422 89004
rect 358630 88952 358636 89004
rect 358688 88992 358694 89004
rect 415394 88992 415400 89004
rect 358688 88964 415400 88992
rect 358688 88952 358694 88964
rect 415394 88952 415400 88964
rect 415452 88952 415458 89004
rect 340414 88680 340420 88732
rect 340472 88720 340478 88732
rect 342530 88720 342536 88732
rect 340472 88692 342536 88720
rect 340472 88680 340478 88692
rect 342530 88680 342536 88692
rect 342588 88680 342594 88732
rect 291838 88272 291844 88324
rect 291896 88312 291902 88324
rect 298002 88312 298008 88324
rect 291896 88284 298008 88312
rect 291896 88272 291902 88284
rect 298002 88272 298008 88284
rect 298060 88272 298066 88324
rect 223482 87592 223488 87644
rect 223540 87632 223546 87644
rect 287698 87632 287704 87644
rect 223540 87604 287704 87632
rect 223540 87592 223546 87604
rect 287698 87592 287704 87604
rect 287756 87592 287762 87644
rect 358814 86912 358820 86964
rect 358872 86952 358878 86964
rect 580166 86952 580172 86964
rect 358872 86924 580172 86952
rect 358872 86912 358878 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 14458 85524 14464 85536
rect 3200 85496 14464 85524
rect 3200 85484 3206 85496
rect 14458 85484 14464 85496
rect 14516 85484 14522 85536
rect 266998 85484 267004 85536
rect 267056 85524 267062 85536
rect 297542 85524 297548 85536
rect 267056 85496 297548 85524
rect 267056 85484 267062 85496
rect 297542 85484 297548 85496
rect 297600 85484 297606 85536
rect 269758 84124 269764 84176
rect 269816 84164 269822 84176
rect 297910 84164 297916 84176
rect 269816 84136 297916 84164
rect 269816 84124 269822 84136
rect 297910 84124 297916 84136
rect 297968 84124 297974 84176
rect 275278 82764 275284 82816
rect 275336 82804 275342 82816
rect 297910 82804 297916 82816
rect 275336 82776 297916 82804
rect 275336 82764 275342 82776
rect 297910 82764 297916 82776
rect 297968 82764 297974 82816
rect 223482 81336 223488 81388
rect 223540 81376 223546 81388
rect 228358 81376 228364 81388
rect 223540 81348 228364 81376
rect 223540 81336 223546 81348
rect 228358 81336 228364 81348
rect 228416 81336 228422 81388
rect 273898 79976 273904 80028
rect 273956 80016 273962 80028
rect 298002 80016 298008 80028
rect 273956 79988 298008 80016
rect 273956 79976 273962 79988
rect 298002 79976 298008 79988
rect 298060 79976 298066 80028
rect 271138 78616 271144 78668
rect 271196 78656 271202 78668
rect 297542 78656 297548 78668
rect 271196 78628 297548 78656
rect 271196 78616 271202 78628
rect 297542 78616 297548 78628
rect 297600 78616 297606 78668
rect 222470 78548 222476 78600
rect 222528 78588 222534 78600
rect 225598 78588 225604 78600
rect 222528 78560 225604 78588
rect 222528 78548 222534 78560
rect 225598 78548 225604 78560
rect 225656 78548 225662 78600
rect 260098 77188 260104 77240
rect 260156 77228 260162 77240
rect 297174 77228 297180 77240
rect 260156 77200 297180 77228
rect 260156 77188 260162 77200
rect 297174 77188 297180 77200
rect 297232 77188 297238 77240
rect 255958 75828 255964 75880
rect 256016 75868 256022 75880
rect 298002 75868 298008 75880
rect 256016 75840 298008 75868
rect 256016 75828 256022 75840
rect 298002 75828 298008 75840
rect 298060 75828 298066 75880
rect 222194 75692 222200 75744
rect 222252 75732 222258 75744
rect 224310 75732 224316 75744
rect 222252 75704 224316 75732
rect 222252 75692 222258 75704
rect 224310 75692 224316 75704
rect 224368 75692 224374 75744
rect 261478 74468 261484 74520
rect 261536 74508 261542 74520
rect 298002 74508 298008 74520
rect 261536 74480 298008 74508
rect 261536 74468 261542 74480
rect 298002 74468 298008 74480
rect 298060 74468 298066 74520
rect 256050 73108 256056 73160
rect 256108 73148 256114 73160
rect 296806 73148 296812 73160
rect 256108 73120 296812 73148
rect 256108 73108 256114 73120
rect 296806 73108 296812 73120
rect 296864 73108 296870 73160
rect 480990 73108 480996 73160
rect 481048 73148 481054 73160
rect 580166 73148 580172 73160
rect 481048 73120 580172 73148
rect 481048 73108 481054 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 222194 73040 222200 73092
rect 222252 73080 222258 73092
rect 224218 73080 224224 73092
rect 222252 73052 224224 73080
rect 222252 73040 222258 73052
rect 224218 73040 224224 73052
rect 224276 73040 224282 73092
rect 223482 70320 223488 70372
rect 223540 70360 223546 70372
rect 250438 70360 250444 70372
rect 223540 70332 250444 70360
rect 223540 70320 223546 70332
rect 250438 70320 250444 70332
rect 250496 70320 250502 70372
rect 265618 70320 265624 70372
rect 265676 70360 265682 70372
rect 298002 70360 298008 70372
rect 265676 70332 298008 70360
rect 265676 70320 265682 70332
rect 298002 70320 298008 70332
rect 298060 70320 298066 70372
rect 343082 69028 343088 69080
rect 343140 69068 343146 69080
rect 489914 69068 489920 69080
rect 343140 69040 489920 69068
rect 343140 69028 343146 69040
rect 489914 69028 489920 69040
rect 489972 69028 489978 69080
rect 268378 68960 268384 69012
rect 268436 69000 268442 69012
rect 297174 69000 297180 69012
rect 268436 68972 297180 69000
rect 268436 68960 268442 68972
rect 297174 68960 297180 68972
rect 297232 68960 297238 69012
rect 223482 67532 223488 67584
rect 223540 67572 223546 67584
rect 235258 67572 235264 67584
rect 223540 67544 235264 67572
rect 223540 67532 223546 67544
rect 235258 67532 235264 67544
rect 235316 67532 235322 67584
rect 282178 67532 282184 67584
rect 282236 67572 282242 67584
rect 297542 67572 297548 67584
rect 282236 67544 297548 67572
rect 282236 67532 282242 67544
rect 297542 67532 297548 67544
rect 297600 67532 297606 67584
rect 343174 66240 343180 66292
rect 343232 66280 343238 66292
rect 482370 66280 482376 66292
rect 343232 66252 482376 66280
rect 343232 66240 343238 66252
rect 482370 66240 482376 66252
rect 482428 66240 482434 66292
rect 222838 64812 222844 64864
rect 222896 64852 222902 64864
rect 233878 64852 233884 64864
rect 222896 64824 233884 64852
rect 222896 64812 222902 64824
rect 233878 64812 233884 64824
rect 233936 64812 233942 64864
rect 278130 64812 278136 64864
rect 278188 64852 278194 64864
rect 297910 64852 297916 64864
rect 278188 64824 297916 64852
rect 278188 64812 278194 64824
rect 297910 64812 297916 64824
rect 297968 64812 297974 64864
rect 343174 63520 343180 63572
rect 343232 63560 343238 63572
rect 418798 63560 418804 63572
rect 343232 63532 418804 63560
rect 343232 63520 343238 63532
rect 418798 63520 418804 63532
rect 418856 63520 418862 63572
rect 342346 62704 342352 62756
rect 342404 62744 342410 62756
rect 343174 62744 343180 62756
rect 342404 62716 343180 62744
rect 342404 62704 342410 62716
rect 343174 62704 343180 62716
rect 343232 62704 343238 62756
rect 342346 62092 342352 62144
rect 342404 62132 342410 62144
rect 480346 62132 480352 62144
rect 342404 62104 480352 62132
rect 342404 62092 342410 62104
rect 480346 62092 480352 62104
rect 480404 62092 480410 62144
rect 264422 62024 264428 62076
rect 264480 62064 264486 62076
rect 298002 62064 298008 62076
rect 264480 62036 298008 62064
rect 264480 62024 264486 62036
rect 298002 62024 298008 62036
rect 298060 62024 298066 62076
rect 215294 61548 215300 61600
rect 215352 61588 215358 61600
rect 342714 61588 342720 61600
rect 215352 61560 342720 61588
rect 215352 61548 215358 61560
rect 342714 61548 342720 61560
rect 342772 61548 342778 61600
rect 168374 61480 168380 61532
rect 168432 61520 168438 61532
rect 341702 61520 341708 61532
rect 168432 61492 341708 61520
rect 168432 61480 168438 61492
rect 341702 61480 341708 61492
rect 341760 61480 341766 61532
rect 158714 61412 158720 61464
rect 158772 61452 158778 61464
rect 343082 61452 343088 61464
rect 158772 61424 343088 61452
rect 158772 61412 158778 61424
rect 343082 61412 343088 61424
rect 343140 61412 343146 61464
rect 154574 61344 154580 61396
rect 154632 61384 154638 61396
rect 342990 61384 342996 61396
rect 154632 61356 342996 61384
rect 154632 61344 154638 61356
rect 342990 61344 342996 61356
rect 343048 61344 343054 61396
rect 356698 60664 356704 60716
rect 356756 60704 356762 60716
rect 580166 60704 580172 60716
rect 356756 60676 580172 60704
rect 356756 60664 356762 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 296622 60188 296628 60240
rect 296680 60228 296686 60240
rect 303614 60228 303620 60240
rect 296680 60200 303620 60228
rect 296680 60188 296686 60200
rect 303614 60188 303620 60200
rect 303672 60188 303678 60240
rect 295242 60120 295248 60172
rect 295300 60160 295306 60172
rect 310514 60160 310520 60172
rect 295300 60132 310520 60160
rect 295300 60120 295306 60132
rect 310514 60120 310520 60132
rect 310572 60120 310578 60172
rect 314654 60120 314660 60172
rect 314712 60160 314718 60172
rect 352558 60160 352564 60172
rect 314712 60132 352564 60160
rect 314712 60120 314718 60132
rect 352558 60120 352564 60132
rect 352616 60120 352622 60172
rect 211154 60052 211160 60104
rect 211212 60092 211218 60104
rect 342806 60092 342812 60104
rect 211212 60064 342812 60092
rect 211212 60052 211218 60064
rect 342806 60052 342812 60064
rect 342864 60052 342870 60104
rect 193214 59984 193220 60036
rect 193272 60024 193278 60036
rect 341334 60024 341340 60036
rect 193272 59996 341340 60024
rect 193272 59984 193278 59996
rect 341334 59984 341340 59996
rect 341392 59984 341398 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 369118 59344 369124 59356
rect 3108 59316 369124 59344
rect 3108 59304 3114 59316
rect 369118 59304 369124 59316
rect 369176 59304 369182 59356
rect 172514 58692 172520 58744
rect 172572 58732 172578 58744
rect 341610 58732 341616 58744
rect 172572 58704 341616 58732
rect 172572 58692 172578 58704
rect 341610 58692 341616 58704
rect 341668 58692 341674 58744
rect 133874 58624 133880 58676
rect 133932 58664 133938 58676
rect 340506 58664 340512 58676
rect 133932 58636 340512 58664
rect 133932 58624 133938 58636
rect 340506 58624 340512 58636
rect 340564 58624 340570 58676
rect 229094 57332 229100 57384
rect 229152 57372 229158 57384
rect 342438 57372 342444 57384
rect 229152 57344 342444 57372
rect 229152 57332 229158 57344
rect 342438 57332 342444 57344
rect 342496 57332 342502 57384
rect 190454 57264 190460 57316
rect 190512 57304 190518 57316
rect 340322 57304 340328 57316
rect 190512 57276 340328 57304
rect 190512 57264 190518 57276
rect 340322 57264 340328 57276
rect 340380 57264 340386 57316
rect 176654 57196 176660 57248
rect 176712 57236 176718 57248
rect 341518 57236 341524 57248
rect 176712 57208 341524 57236
rect 176712 57196 176718 57208
rect 341518 57196 341524 57208
rect 341576 57196 341582 57248
rect 233234 55972 233240 56024
rect 233292 56012 233298 56024
rect 343174 56012 343180 56024
rect 233292 55984 343180 56012
rect 233292 55972 233298 55984
rect 343174 55972 343180 55984
rect 343232 55972 343238 56024
rect 226334 55904 226340 55956
rect 226392 55944 226398 55956
rect 341242 55944 341248 55956
rect 226392 55916 341248 55944
rect 226392 55904 226398 55916
rect 341242 55904 341248 55916
rect 341300 55904 341306 55956
rect 179414 55836 179420 55888
rect 179472 55876 179478 55888
rect 341426 55876 341432 55888
rect 179472 55848 341432 55876
rect 179472 55836 179478 55848
rect 341426 55836 341432 55848
rect 341484 55836 341490 55888
rect 247034 54612 247040 54664
rect 247092 54652 247098 54664
rect 340138 54652 340144 54664
rect 247092 54624 340144 54652
rect 247092 54612 247098 54624
rect 340138 54612 340144 54624
rect 340196 54612 340202 54664
rect 218054 54544 218060 54596
rect 218112 54584 218118 54596
rect 342622 54584 342628 54596
rect 218112 54556 342628 54584
rect 218112 54544 218118 54556
rect 342622 54544 342628 54556
rect 342680 54544 342686 54596
rect 204254 54476 204260 54528
rect 204312 54516 204318 54528
rect 340230 54516 340236 54528
rect 204312 54488 340236 54516
rect 204312 54476 204318 54488
rect 340230 54476 340236 54488
rect 340288 54476 340294 54528
rect 346394 53048 346400 53100
rect 346452 53088 346458 53100
rect 509786 53088 509792 53100
rect 346452 53060 509792 53088
rect 346452 53048 346458 53060
rect 509786 53048 509792 53060
rect 509844 53048 509850 53100
rect 251174 50328 251180 50380
rect 251232 50368 251238 50380
rect 341058 50368 341064 50380
rect 251232 50340 341064 50368
rect 251232 50328 251238 50340
rect 341058 50328 341064 50340
rect 341116 50328 341122 50380
rect 201494 47540 201500 47592
rect 201552 47580 201558 47592
rect 491938 47580 491944 47592
rect 201552 47552 491944 47580
rect 201552 47540 201558 47552
rect 491938 47540 491944 47552
rect 491996 47540 492002 47592
rect 359550 46860 359556 46912
rect 359608 46900 359614 46912
rect 580166 46900 580172 46912
rect 359608 46872 580172 46900
rect 359608 46860 359614 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 472710 45540 472716 45552
rect 3476 45512 472716 45540
rect 3476 45500 3482 45512
rect 472710 45500 472716 45512
rect 472768 45500 472774 45552
rect 99374 43392 99380 43444
rect 99432 43432 99438 43444
rect 513006 43432 513012 43444
rect 99432 43404 513012 43432
rect 99432 43392 99438 43404
rect 513006 43392 513012 43404
rect 513064 43392 513070 43444
rect 151814 42032 151820 42084
rect 151872 42072 151878 42084
rect 342898 42072 342904 42084
rect 151872 42044 342904 42072
rect 151872 42032 151878 42044
rect 342898 42032 342904 42044
rect 342956 42032 342962 42084
rect 208394 40808 208400 40860
rect 208452 40848 208458 40860
rect 341150 40848 341156 40860
rect 208452 40820 341156 40848
rect 208452 40808 208458 40820
rect 341150 40808 341156 40820
rect 341208 40808 341214 40860
rect 120074 40740 120080 40792
rect 120132 40780 120138 40792
rect 481266 40780 481272 40792
rect 120132 40752 481272 40780
rect 120132 40740 120138 40752
rect 481266 40740 481272 40752
rect 481324 40740 481330 40792
rect 56594 40672 56600 40724
rect 56652 40712 56658 40724
rect 512270 40712 512276 40724
rect 56652 40684 512276 40712
rect 56652 40672 56658 40684
rect 512270 40672 512276 40684
rect 512328 40672 512334 40724
rect 113174 37884 113180 37936
rect 113232 37924 113238 37936
rect 462958 37924 462964 37936
rect 113232 37896 462964 37924
rect 113232 37884 113238 37896
rect 462958 37884 462964 37896
rect 463016 37884 463022 37936
rect 117314 36524 117320 36576
rect 117372 36564 117378 36576
rect 436738 36564 436744 36576
rect 117372 36536 436744 36564
rect 117372 36524 117378 36536
rect 436738 36524 436744 36536
rect 436796 36524 436802 36576
rect 235994 35300 236000 35352
rect 236052 35340 236058 35352
rect 340046 35340 340052 35352
rect 236052 35312 340052 35340
rect 236052 35300 236058 35312
rect 340046 35300 340052 35312
rect 340104 35300 340110 35352
rect 110414 35232 110420 35284
rect 110472 35272 110478 35284
rect 496170 35272 496176 35284
rect 110472 35244 496176 35272
rect 110472 35232 110478 35244
rect 496170 35232 496176 35244
rect 496228 35232 496234 35284
rect 23474 35164 23480 35216
rect 23532 35204 23538 35216
rect 416038 35204 416044 35216
rect 23532 35176 416044 35204
rect 23532 35164 23538 35176
rect 416038 35164 416044 35176
rect 416096 35164 416102 35216
rect 70394 33736 70400 33788
rect 70452 33776 70458 33788
rect 501230 33776 501236 33788
rect 70452 33748 501236 33776
rect 70452 33736 70458 33748
rect 501230 33736 501236 33748
rect 501288 33736 501294 33788
rect 480898 33056 480904 33108
rect 480956 33096 480962 33108
rect 580166 33096 580172 33108
rect 480956 33068 580172 33096
rect 480956 33056 480962 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 378134 31016 378140 31068
rect 378192 31056 378198 31068
rect 476850 31056 476856 31068
rect 378192 31028 476856 31056
rect 378192 31016 378198 31028
rect 476850 31016 476856 31028
rect 476908 31016 476914 31068
rect 77294 29588 77300 29640
rect 77352 29628 77358 29640
rect 502978 29628 502984 29640
rect 77352 29600 502984 29628
rect 77352 29588 77358 29600
rect 502978 29588 502984 29600
rect 503036 29588 503042 29640
rect 92474 26868 92480 26920
rect 92532 26908 92538 26920
rect 493410 26908 493416 26920
rect 92532 26880 493416 26908
rect 92532 26868 92538 26880
rect 493410 26868 493416 26880
rect 493468 26868 493474 26920
rect 371234 22720 371240 22772
rect 371292 22760 371298 22772
rect 440878 22760 440884 22772
rect 371292 22732 440884 22760
rect 371292 22720 371298 22732
rect 440878 22720 440884 22732
rect 440936 22720 440942 22772
rect 396166 21428 396172 21480
rect 396224 21468 396230 21480
rect 422938 21468 422944 21480
rect 396224 21440 422944 21468
rect 396224 21428 396230 21440
rect 422938 21428 422944 21440
rect 422996 21428 423002 21480
rect 423766 21428 423772 21480
rect 423824 21468 423830 21480
rect 504450 21468 504456 21480
rect 423824 21440 504456 21468
rect 423824 21428 423830 21440
rect 504450 21428 504456 21440
rect 504508 21428 504514 21480
rect 60734 21360 60740 21412
rect 60792 21400 60798 21412
rect 475470 21400 475476 21412
rect 60792 21372 475476 21400
rect 60792 21360 60798 21372
rect 475470 21360 475476 21372
rect 475528 21360 475534 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 510706 20652 510712 20664
rect 3476 20624 510712 20652
rect 3476 20612 3482 20624
rect 510706 20612 510712 20624
rect 510764 20612 510770 20664
rect 102134 19932 102140 19984
rect 102192 19972 102198 19984
rect 496078 19972 496084 19984
rect 102192 19944 496084 19972
rect 102192 19932 102198 19944
rect 496078 19932 496084 19944
rect 496136 19932 496142 19984
rect 197354 18708 197360 18760
rect 197412 18748 197418 18760
rect 340966 18748 340972 18760
rect 197412 18720 340972 18748
rect 197412 18708 197418 18720
rect 340966 18708 340972 18720
rect 341024 18708 341030 18760
rect 360194 18708 360200 18760
rect 360252 18748 360258 18760
rect 450538 18748 450544 18760
rect 360252 18720 450544 18748
rect 360252 18708 360258 18720
rect 450538 18708 450544 18720
rect 450596 18708 450602 18760
rect 106274 18640 106280 18692
rect 106332 18680 106338 18692
rect 404998 18680 405004 18692
rect 106332 18652 405004 18680
rect 106332 18640 106338 18652
rect 404998 18640 405004 18652
rect 405056 18640 405062 18692
rect 19334 18572 19340 18624
rect 19392 18612 19398 18624
rect 402238 18612 402244 18624
rect 19392 18584 402244 18612
rect 19392 18572 19398 18584
rect 402238 18572 402244 18584
rect 402296 18572 402302 18624
rect 420178 17280 420184 17332
rect 420236 17320 420242 17332
rect 498286 17320 498292 17332
rect 420236 17292 498292 17320
rect 420236 17280 420242 17292
rect 498286 17280 498292 17292
rect 498344 17280 498350 17332
rect 357434 17212 357440 17264
rect 357492 17252 357498 17264
rect 454678 17252 454684 17264
rect 357492 17224 454684 17252
rect 357492 17212 357498 17224
rect 454678 17212 454684 17224
rect 454736 17212 454742 17264
rect 390922 15920 390928 15972
rect 390980 15960 390986 15972
rect 440234 15960 440240 15972
rect 390980 15932 440240 15960
rect 390980 15920 390986 15932
rect 440234 15920 440240 15932
rect 440292 15920 440298 15972
rect 81618 15852 81624 15904
rect 81676 15892 81682 15904
rect 493318 15892 493324 15904
rect 81676 15864 493324 15892
rect 81676 15852 81682 15864
rect 493318 15852 493324 15864
rect 493376 15852 493382 15904
rect 254210 14424 254216 14476
rect 254268 14464 254274 14476
rect 494790 14464 494796 14476
rect 254268 14436 494796 14464
rect 254268 14424 254274 14436
rect 494790 14424 494796 14436
rect 494848 14424 494854 14476
rect 353570 13064 353576 13116
rect 353628 13104 353634 13116
rect 476758 13104 476764 13116
rect 353628 13076 476764 13104
rect 353628 13064 353634 13076
rect 476758 13064 476764 13076
rect 476816 13064 476822 13116
rect 378686 11704 378692 11756
rect 378744 11744 378750 11756
rect 455690 11744 455696 11756
rect 378744 11716 455696 11744
rect 378744 11704 378750 11716
rect 455690 11704 455696 11716
rect 455748 11704 455754 11756
rect 242894 10344 242900 10396
rect 242952 10384 242958 10396
rect 342254 10384 342260 10396
rect 242952 10356 342260 10384
rect 242952 10344 242958 10356
rect 342254 10344 342260 10356
rect 342312 10344 342318 10396
rect 240134 10276 240140 10328
rect 240192 10316 240198 10328
rect 340874 10316 340880 10328
rect 240192 10288 340880 10316
rect 240192 10276 240198 10288
rect 340874 10276 340880 10288
rect 340932 10276 340938 10328
rect 477862 10276 477868 10328
rect 477920 10316 477926 10328
rect 494698 10316 494704 10328
rect 477920 10288 494704 10316
rect 477920 10276 477926 10288
rect 494698 10276 494704 10288
rect 494756 10276 494762 10328
rect 445018 9052 445024 9104
rect 445076 9092 445082 9104
rect 494698 9092 494704 9104
rect 445076 9064 494704 9092
rect 445076 9052 445082 9064
rect 494698 9052 494704 9064
rect 494756 9052 494762 9104
rect 89162 8984 89168 9036
rect 89220 9024 89226 9036
rect 510338 9024 510344 9036
rect 89220 8996 510344 9024
rect 89220 8984 89226 8996
rect 510338 8984 510344 8996
rect 510396 8984 510402 9036
rect 85666 8916 85672 8968
rect 85724 8956 85730 8968
rect 509970 8956 509976 8968
rect 85724 8928 509976 8956
rect 85724 8916 85730 8928
rect 509970 8916 509976 8928
rect 510028 8916 510034 8968
rect 396074 8236 396080 8288
rect 396132 8276 396138 8288
rect 402514 8276 402520 8288
rect 396132 8248 402520 8276
rect 396132 8236 396138 8248
rect 402514 8236 402520 8248
rect 402572 8236 402578 8288
rect 482370 8236 482376 8288
rect 482428 8276 482434 8288
rect 487614 8276 487620 8288
rect 482428 8248 487620 8276
rect 482428 8236 482434 8248
rect 487614 8236 487620 8248
rect 487672 8236 487678 8288
rect 418798 7760 418804 7812
rect 418856 7800 418862 7812
rect 484026 7800 484032 7812
rect 418856 7772 484032 7800
rect 418856 7760 418862 7772
rect 484026 7760 484032 7772
rect 484084 7760 484090 7812
rect 67910 7692 67916 7744
rect 67968 7732 67974 7744
rect 475378 7732 475384 7744
rect 67968 7704 475384 7732
rect 67968 7692 67974 7704
rect 475378 7692 475384 7704
rect 475436 7692 475442 7744
rect 478690 7692 478696 7744
rect 478748 7732 478754 7744
rect 580994 7732 581000 7744
rect 478748 7704 581000 7732
rect 478748 7692 478754 7704
rect 580994 7692 581000 7704
rect 581052 7692 581058 7744
rect 64322 7624 64328 7676
rect 64380 7664 64386 7676
rect 512822 7664 512828 7676
rect 64380 7636 512828 7664
rect 64380 7624 64386 7636
rect 512822 7624 512828 7636
rect 512880 7624 512886 7676
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 510614 7596 510620 7608
rect 4120 7568 510620 7596
rect 4120 7556 4126 7568
rect 510614 7556 510620 7568
rect 510672 7556 510678 7608
rect 359458 6808 359464 6860
rect 359516 6848 359522 6860
rect 580166 6848 580172 6860
rect 359516 6820 580172 6848
rect 359516 6808 359522 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 46658 6264 46664 6316
rect 46716 6304 46722 6316
rect 489638 6304 489644 6316
rect 46716 6276 489644 6304
rect 46716 6264 46722 6276
rect 489638 6264 489644 6276
rect 489696 6264 489702 6316
rect 35986 6196 35992 6248
rect 36044 6236 36050 6248
rect 491570 6236 491576 6248
rect 36044 6208 491576 6236
rect 36044 6196 36050 6208
rect 491570 6196 491576 6208
rect 491628 6196 491634 6248
rect 39574 6128 39580 6180
rect 39632 6168 39638 6180
rect 499942 6168 499948 6180
rect 39632 6140 499948 6168
rect 39632 6128 39638 6140
rect 499942 6128 499948 6140
rect 500000 6128 500006 6180
rect 141234 4972 141240 5024
rect 141292 5012 141298 5024
rect 141292 4984 142154 5012
rect 141292 4972 141298 4984
rect 142126 4944 142154 4984
rect 357618 4972 357624 5024
rect 357676 5012 357682 5024
rect 473446 5012 473452 5024
rect 357676 4984 473452 5012
rect 357676 4972 357682 4984
rect 473446 4972 473452 4984
rect 473504 4972 473510 5024
rect 477954 4972 477960 5024
rect 478012 5012 478018 5024
rect 559742 5012 559748 5024
rect 478012 4984 559748 5012
rect 478012 4972 478018 4984
rect 559742 4972 559748 4984
rect 559800 4972 559806 5024
rect 342530 4944 342536 4956
rect 142126 4916 342536 4944
rect 342530 4904 342536 4916
rect 342588 4904 342594 4956
rect 350442 4904 350448 4956
rect 350500 4944 350506 4956
rect 508314 4944 508320 4956
rect 350500 4916 508320 4944
rect 350500 4904 350506 4916
rect 508314 4904 508320 4916
rect 508372 4904 508378 4956
rect 50154 4836 50160 4888
rect 50212 4876 50218 4888
rect 507670 4876 507676 4888
rect 50212 4848 507676 4876
rect 50212 4836 50218 4848
rect 507670 4836 507676 4848
rect 507728 4836 507734 4888
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 512730 4808 512736 4820
rect 2924 4780 512736 4808
rect 2924 4768 2930 4780
rect 512730 4768 512736 4780
rect 512788 4768 512794 4820
rect 339862 3952 339868 4004
rect 339920 3992 339926 4004
rect 353386 3992 353392 4004
rect 339920 3964 353392 3992
rect 339920 3952 339926 3964
rect 353386 3952 353392 3964
rect 353444 3952 353450 4004
rect 332686 3884 332692 3936
rect 332744 3924 332750 3936
rect 350534 3924 350540 3936
rect 332744 3896 350540 3924
rect 332744 3884 332750 3896
rect 350534 3884 350540 3896
rect 350592 3884 350598 3936
rect 336274 3816 336280 3868
rect 336332 3856 336338 3868
rect 355410 3856 355416 3868
rect 336332 3828 355416 3856
rect 336332 3816 336338 3828
rect 355410 3816 355416 3828
rect 355468 3816 355474 3868
rect 296530 3748 296536 3800
rect 296588 3788 296594 3800
rect 322106 3788 322112 3800
rect 296588 3760 322112 3788
rect 296588 3748 296594 3760
rect 322106 3748 322112 3760
rect 322164 3748 322170 3800
rect 325602 3748 325608 3800
rect 325660 3788 325666 3800
rect 351178 3788 351184 3800
rect 325660 3760 351184 3788
rect 325660 3748 325666 3760
rect 351178 3748 351184 3760
rect 351236 3748 351242 3800
rect 307938 3680 307944 3732
rect 307996 3720 308002 3732
rect 355318 3720 355324 3732
rect 307996 3692 355324 3720
rect 307996 3680 308002 3692
rect 355318 3680 355324 3692
rect 355376 3680 355382 3732
rect 538858 3680 538864 3732
rect 538916 3720 538922 3732
rect 556154 3720 556160 3732
rect 538916 3692 556160 3720
rect 538916 3680 538922 3692
rect 556154 3680 556160 3692
rect 556212 3680 556218 3732
rect 222746 3612 222752 3664
rect 222804 3652 222810 3664
rect 340414 3652 340420 3664
rect 222804 3624 340420 3652
rect 222804 3612 222810 3624
rect 340414 3612 340420 3624
rect 340472 3612 340478 3664
rect 343358 3612 343364 3664
rect 343416 3652 343422 3664
rect 353294 3652 353300 3664
rect 343416 3624 353300 3652
rect 343416 3612 343422 3624
rect 353294 3612 353300 3624
rect 353352 3612 353358 3664
rect 453298 3612 453304 3664
rect 453356 3652 453362 3664
rect 508498 3652 508504 3664
rect 453356 3624 508504 3652
rect 453356 3612 453362 3624
rect 508498 3612 508504 3624
rect 508556 3612 508562 3664
rect 530578 3612 530584 3664
rect 530636 3652 530642 3664
rect 530636 3624 531452 3652
rect 530636 3612 530642 3624
rect 102134 3544 102140 3596
rect 102192 3584 102198 3596
rect 103330 3584 103336 3596
rect 102192 3556 103336 3584
rect 102192 3544 102198 3556
rect 103330 3544 103336 3556
rect 103388 3544 103394 3596
rect 124674 3544 124680 3596
rect 124732 3584 124738 3596
rect 488994 3584 489000 3596
rect 124732 3556 489000 3584
rect 124732 3544 124738 3556
rect 488994 3544 489000 3556
rect 489052 3544 489058 3596
rect 526438 3544 526444 3596
rect 526496 3584 526502 3596
rect 531314 3584 531320 3596
rect 526496 3556 531320 3584
rect 526496 3544 526502 3556
rect 531314 3544 531320 3556
rect 531372 3544 531378 3596
rect 531424 3584 531452 3624
rect 531958 3612 531964 3664
rect 532016 3652 532022 3664
rect 541986 3652 541992 3664
rect 532016 3624 541992 3652
rect 532016 3612 532022 3624
rect 541986 3612 541992 3624
rect 542044 3612 542050 3664
rect 538398 3584 538404 3596
rect 531424 3556 538404 3584
rect 538398 3544 538404 3556
rect 538456 3544 538462 3596
rect 544378 3544 544384 3596
rect 544436 3584 544442 3596
rect 573910 3584 573916 3596
rect 544436 3556 573916 3584
rect 544436 3544 544442 3556
rect 573910 3544 573916 3556
rect 573968 3544 573974 3596
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 472618 3516 472624 3528
rect 32456 3488 472624 3516
rect 32456 3476 32462 3488
rect 472618 3476 472624 3488
rect 472676 3476 472682 3528
rect 479426 3476 479432 3528
rect 479484 3516 479490 3528
rect 485222 3516 485228 3528
rect 479484 3488 485228 3516
rect 479484 3476 479490 3488
rect 485222 3476 485228 3488
rect 485280 3476 485286 3528
rect 498194 3476 498200 3528
rect 498252 3516 498258 3528
rect 499022 3516 499028 3528
rect 498252 3488 499028 3516
rect 498252 3476 498258 3488
rect 499022 3476 499028 3488
rect 499080 3476 499086 3528
rect 522298 3476 522304 3528
rect 522356 3516 522362 3528
rect 524230 3516 524236 3528
rect 522356 3488 524236 3516
rect 522356 3476 522362 3488
rect 524230 3476 524236 3488
rect 524288 3476 524294 3528
rect 525058 3476 525064 3528
rect 525116 3516 525122 3528
rect 527818 3516 527824 3528
rect 525116 3488 527824 3516
rect 525116 3476 525122 3488
rect 527818 3476 527824 3488
rect 527876 3476 527882 3528
rect 534718 3476 534724 3528
rect 534776 3516 534782 3528
rect 534776 3488 538214 3516
rect 534776 3476 534782 3488
rect 28902 3408 28908 3460
rect 28960 3448 28966 3460
rect 468478 3448 468484 3460
rect 28960 3420 468484 3448
rect 28960 3408 28966 3420
rect 468478 3408 468484 3420
rect 468536 3408 468542 3460
rect 482278 3408 482284 3460
rect 482336 3448 482342 3460
rect 510062 3448 510068 3460
rect 482336 3420 510068 3448
rect 482336 3408 482342 3420
rect 510062 3408 510068 3420
rect 510120 3408 510126 3460
rect 527910 3408 527916 3460
rect 527968 3448 527974 3460
rect 534902 3448 534908 3460
rect 527968 3420 534908 3448
rect 527968 3408 527974 3420
rect 534902 3408 534908 3420
rect 534960 3408 534966 3460
rect 538186 3448 538214 3488
rect 549898 3476 549904 3528
rect 549956 3516 549962 3528
rect 549956 3488 578832 3516
rect 549956 3476 549962 3488
rect 545482 3448 545488 3460
rect 538186 3420 545488 3448
rect 545482 3408 545488 3420
rect 545540 3408 545546 3460
rect 545758 3408 545764 3460
rect 545816 3448 545822 3460
rect 577406 3448 577412 3460
rect 545816 3420 577412 3448
rect 545816 3408 545822 3420
rect 577406 3408 577412 3420
rect 577464 3408 577470 3460
rect 578804 3448 578832 3488
rect 578878 3476 578884 3528
rect 578936 3516 578942 3528
rect 579798 3516 579804 3528
rect 578936 3488 579804 3516
rect 578936 3476 578942 3488
rect 579798 3476 579804 3488
rect 579856 3476 579862 3528
rect 582190 3448 582196 3460
rect 578804 3420 582196 3448
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 143534 3340 143540 3392
rect 143592 3380 143598 3392
rect 144730 3380 144736 3392
rect 143592 3352 144736 3380
rect 143592 3340 143598 3352
rect 144730 3340 144736 3352
rect 144788 3340 144794 3392
rect 168374 3340 168380 3392
rect 168432 3380 168438 3392
rect 169570 3380 169576 3392
rect 168432 3352 169576 3380
rect 168432 3340 168438 3352
rect 169570 3340 169576 3352
rect 169628 3340 169634 3392
rect 193214 3340 193220 3392
rect 193272 3380 193278 3392
rect 194410 3380 194416 3392
rect 193272 3352 194416 3380
rect 193272 3340 193278 3352
rect 194410 3340 194416 3352
rect 194468 3340 194474 3392
rect 218054 3340 218060 3392
rect 218112 3380 218118 3392
rect 219250 3380 219256 3392
rect 218112 3352 219256 3380
rect 218112 3340 218118 3352
rect 219250 3340 219256 3352
rect 219308 3340 219314 3392
rect 242894 3340 242900 3392
rect 242952 3380 242958 3392
rect 244090 3380 244096 3392
rect 242952 3352 244096 3380
rect 242952 3340 242958 3352
rect 244090 3340 244096 3352
rect 244148 3340 244154 3392
rect 414658 3340 414664 3392
rect 414716 3380 414722 3392
rect 420178 3380 420184 3392
rect 414716 3352 420184 3380
rect 414716 3340 414722 3352
rect 420178 3340 420184 3352
rect 420236 3340 420242 3392
rect 423766 3340 423772 3392
rect 423824 3380 423830 3392
rect 424962 3380 424968 3392
rect 423824 3352 424968 3380
rect 423824 3340 423830 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 448514 3340 448520 3392
rect 448572 3380 448578 3392
rect 449802 3380 449808 3392
rect 448572 3352 449808 3380
rect 448572 3340 448578 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 398834 3136 398840 3188
rect 398892 3176 398898 3188
rect 400122 3176 400128 3188
rect 398892 3148 400128 3176
rect 398892 3136 398898 3148
rect 400122 3136 400128 3148
rect 400180 3136 400186 3188
rect 415394 3136 415400 3188
rect 415452 3176 415458 3188
rect 416682 3176 416688 3188
rect 415452 3148 416688 3176
rect 415452 3136 415458 3148
rect 416682 3136 416688 3148
rect 416740 3136 416746 3188
rect 440234 3136 440240 3188
rect 440292 3176 440298 3188
rect 441522 3176 441528 3188
rect 440292 3148 441528 3176
rect 440292 3136 440298 3148
rect 441522 3136 441528 3148
rect 441580 3136 441586 3188
rect 506474 3136 506480 3188
rect 506532 3176 506538 3188
rect 508958 3176 508964 3188
rect 506532 3148 508964 3176
rect 506532 3136 506538 3148
rect 508958 3136 508964 3148
rect 509016 3136 509022 3188
rect 373994 3000 374000 3052
rect 374052 3040 374058 3052
rect 375282 3040 375288 3052
rect 374052 3012 375288 3040
rect 374052 3000 374058 3012
rect 375282 3000 375288 3012
rect 375340 3000 375346 3052
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 235172 700612 235224 700664
rect 253296 700612 253348 700664
rect 218980 700544 219032 700596
rect 253388 700544 253440 700596
rect 154120 700476 154172 700528
rect 264336 700476 264388 700528
rect 283840 700476 283892 700528
rect 477040 700476 477092 700528
rect 89168 700408 89220 700460
rect 265624 700408 265676 700460
rect 300124 700408 300176 700460
rect 320916 700408 320968 700460
rect 360844 700408 360896 700460
rect 559656 700408 559708 700460
rect 72976 700340 73028 700392
rect 253204 700340 253256 700392
rect 317420 700340 317472 700392
rect 543464 700340 543516 700392
rect 24308 700272 24360 700324
rect 406384 700272 406436 700324
rect 520924 699660 520976 699712
rect 527180 699660 527232 699712
rect 397460 698912 397512 698964
rect 477132 698912 477184 698964
rect 266360 697620 266412 697672
rect 267648 697620 267700 697672
rect 105452 697552 105504 697604
rect 337384 697552 337436 697604
rect 525156 696940 525208 696992
rect 580172 696940 580224 696992
rect 316132 683136 316184 683188
rect 580172 683136 580224 683188
rect 403716 670692 403768 670744
rect 580172 670692 580224 670744
rect 6920 665796 6972 665848
rect 475752 665796 475804 665848
rect 52092 663824 52144 663876
rect 355416 663824 355468 663876
rect 46480 663756 46532 663808
rect 352564 663756 352616 663808
rect 50436 663076 50488 663128
rect 279424 663076 279476 663128
rect 46756 663008 46808 663060
rect 279976 663008 280028 663060
rect 51724 662940 51776 662992
rect 352840 662940 352892 662992
rect 51080 662872 51132 662924
rect 352656 662872 352708 662924
rect 50896 662804 50948 662856
rect 353024 662804 353076 662856
rect 52000 662736 52052 662788
rect 355324 662736 355376 662788
rect 47860 662668 47912 662720
rect 352932 662668 352984 662720
rect 45468 662600 45520 662652
rect 352748 662600 352800 662652
rect 51908 662532 51960 662584
rect 405096 662532 405148 662584
rect 52184 662464 52236 662516
rect 405740 662464 405792 662516
rect 46388 662396 46440 662448
rect 403808 662396 403860 662448
rect 201500 661784 201552 661836
rect 422944 661784 422996 661836
rect 50252 661716 50304 661768
rect 279332 661716 279384 661768
rect 136640 661648 136692 661700
rect 475660 661648 475712 661700
rect 50528 661580 50580 661632
rect 280068 661580 280120 661632
rect 49148 661512 49200 661564
rect 279516 661512 279568 661564
rect 50804 661444 50856 661496
rect 356888 661444 356940 661496
rect 50620 661376 50672 661428
rect 401600 661376 401652 661428
rect 51816 661308 51868 661360
rect 405832 661308 405884 661360
rect 49792 661240 49844 661292
rect 512000 661240 512052 661292
rect 3608 661172 3660 661224
rect 478880 661172 478932 661224
rect 3424 661104 3476 661156
rect 484400 661104 484452 661156
rect 3792 661036 3844 661088
rect 498200 661036 498252 661088
rect 49424 660560 49476 660612
rect 257436 660560 257488 660612
rect 49608 660492 49660 660544
rect 278136 660492 278188 660544
rect 50160 660424 50212 660476
rect 488540 660424 488592 660476
rect 50712 660356 50764 660408
rect 279608 660356 279660 660408
rect 50344 660288 50396 660340
rect 500960 660288 501012 660340
rect 49516 660220 49568 660272
rect 279056 660220 279108 660272
rect 49240 660152 49292 660204
rect 279148 660152 279200 660204
rect 48228 660084 48280 660136
rect 278964 660084 279016 660136
rect 46848 660016 46900 660068
rect 279240 660016 279292 660068
rect 51356 659948 51408 660000
rect 296904 659948 296956 660000
rect 51264 659880 51316 659932
rect 356980 659880 357032 659932
rect 3332 659812 3384 659864
rect 477224 659812 477276 659864
rect 50344 658656 50396 658708
rect 50988 658656 51040 658708
rect 254584 656888 254636 656940
rect 353116 656888 353168 656940
rect 48688 652740 48740 652792
rect 49976 652740 50028 652792
rect 50988 651380 51040 651432
rect 52184 651380 52236 651432
rect 49240 648524 49292 648576
rect 50160 648524 50212 648576
rect 253940 645872 253992 645924
rect 257344 645872 257396 645924
rect 526444 643084 526496 643136
rect 580172 643084 580224 643136
rect 357348 642812 357400 642864
rect 371700 642812 371752 642864
rect 361028 642744 361080 642796
rect 379980 642744 380032 642796
rect 353208 642676 353260 642728
rect 382188 642676 382240 642728
rect 357256 642608 357308 642660
rect 388812 642608 388864 642660
rect 392676 642608 392728 642660
rect 399300 642608 399352 642660
rect 359464 642540 359516 642592
rect 376116 642540 376168 642592
rect 376208 642540 376260 642592
rect 400312 642540 400364 642592
rect 370044 642472 370096 642524
rect 403164 642472 403216 642524
rect 310428 642404 310480 642456
rect 361764 642404 361816 642456
rect 366180 642404 366232 642456
rect 399116 642404 399168 642456
rect 287612 642336 287664 642388
rect 351368 642336 351420 642388
rect 355968 642336 356020 642388
rect 391020 642336 391072 642388
rect 392124 642336 392176 642388
rect 399208 642336 399260 642388
rect 293132 642268 293184 642320
rect 321100 642268 321152 642320
rect 365536 642268 365588 642320
rect 383292 642268 383344 642320
rect 393228 642268 393280 642320
rect 400496 642268 400548 642320
rect 295248 642200 295300 642252
rect 323676 642200 323728 642252
rect 349896 642200 349948 642252
rect 377772 642200 377824 642252
rect 387156 642200 387208 642252
rect 400956 642200 401008 642252
rect 300768 642132 300820 642184
rect 329196 642132 329248 642184
rect 355600 642132 355652 642184
rect 386052 642132 386104 642184
rect 394332 642132 394384 642184
rect 405280 642132 405332 642184
rect 286508 642064 286560 642116
rect 321008 642064 321060 642116
rect 371148 642064 371200 642116
rect 399668 642064 399720 642116
rect 296352 641996 296404 642048
rect 331864 641996 331916 642048
rect 333244 641996 333296 642048
rect 363420 641996 363472 642048
rect 374460 641996 374512 642048
rect 405188 641996 405240 642048
rect 284208 641928 284260 641980
rect 325056 641928 325108 641980
rect 359740 641928 359792 641980
rect 373356 641928 373408 641980
rect 290924 641860 290976 641912
rect 319444 641860 319496 641912
rect 357072 641860 357124 641912
rect 381084 641860 381136 641912
rect 394884 641860 394936 641912
rect 400588 641860 400640 641912
rect 297548 641792 297600 641844
rect 349804 641792 349856 641844
rect 360108 641792 360160 641844
rect 368388 641792 368440 641844
rect 378048 641792 378100 641844
rect 386604 641792 386656 641844
rect 393780 641792 393832 641844
rect 399392 641792 399444 641844
rect 472624 641792 472676 641844
rect 493232 641792 493284 641844
rect 49056 641724 49108 641776
rect 50252 641724 50304 641776
rect 358820 641724 358872 641776
rect 366732 641724 366784 641776
rect 375564 641724 375616 641776
rect 376208 641724 376260 641776
rect 395436 641724 395488 641776
rect 399760 641724 399812 641776
rect 405004 641724 405056 641776
rect 510620 641724 510672 641776
rect 358544 641180 358596 641232
rect 391572 641180 391624 641232
rect 278688 641112 278740 641164
rect 398472 641112 398524 641164
rect 315856 641044 315908 641096
rect 523684 641044 523736 641096
rect 278596 640976 278648 641028
rect 310428 640976 310480 641028
rect 314108 640976 314160 641028
rect 530584 640976 530636 641028
rect 355508 640908 355560 640960
rect 378324 640908 378376 640960
rect 357164 640840 357216 640892
rect 383844 640840 383896 640892
rect 357808 640772 357860 640824
rect 388260 640772 388312 640824
rect 359188 640704 359240 640756
rect 389364 640704 389416 640756
rect 313004 640636 313056 640688
rect 338764 640636 338816 640688
rect 342904 640636 342956 640688
rect 384948 640636 385000 640688
rect 387708 640636 387760 640688
rect 401876 640636 401928 640688
rect 308588 640568 308640 640620
rect 356796 640568 356848 640620
rect 389916 640568 389968 640620
rect 401600 640568 401652 640620
rect 303068 640500 303120 640552
rect 356704 640500 356756 640552
rect 357900 640500 357952 640552
rect 396540 640500 396592 640552
rect 315212 640432 315264 640484
rect 322388 640432 322440 640484
rect 360016 640432 360068 640484
rect 379428 640432 379480 640484
rect 310336 640364 310388 640416
rect 320824 640364 320876 640416
rect 361212 640364 361264 640416
rect 384396 640364 384448 640416
rect 254492 640296 254544 640348
rect 273996 640296 274048 640348
rect 311808 640296 311860 640348
rect 323584 640296 323636 640348
rect 361120 640296 361172 640348
rect 385500 640296 385552 640348
rect 367560 639956 367612 640008
rect 364800 639888 364852 639940
rect 373264 639888 373316 639940
rect 365720 639820 365772 639872
rect 373172 639820 373224 639872
rect 368112 639752 368164 639804
rect 372344 639752 372396 639804
rect 327724 639684 327776 639736
rect 382372 639684 382424 639736
rect 358452 639616 358504 639668
rect 374644 639616 374696 639668
rect 377496 639616 377548 639668
rect 358636 639548 358688 639600
rect 376300 639548 376352 639600
rect 319720 639480 319772 639532
rect 378508 639480 378560 639532
rect 319536 639412 319588 639464
rect 380164 639412 380216 639464
rect 319168 639344 319220 639396
rect 322480 639344 322532 639396
rect 358912 639344 358964 639396
rect 371884 639344 371936 639396
rect 372344 639344 372396 639396
rect 373080 639344 373132 639396
rect 373172 639344 373224 639396
rect 373264 639344 373316 639396
rect 374000 639344 374052 639396
rect 292028 639276 292080 639328
rect 294052 639276 294104 639328
rect 305092 639276 305144 639328
rect 307484 639276 307536 639328
rect 309692 639276 309744 639328
rect 354036 639276 354088 639328
rect 370596 639276 370648 639328
rect 351276 639208 351328 639260
rect 353944 639140 353996 639192
rect 322204 639072 322256 639124
rect 361488 639004 361540 639056
rect 322296 638936 322348 638988
rect 381268 639344 381320 639396
rect 385684 639548 385736 639600
rect 381728 639344 381780 639396
rect 401784 639548 401836 639600
rect 396264 639412 396316 639464
rect 399024 639412 399076 639464
rect 385868 639344 385920 639396
rect 385960 639344 386012 639396
rect 386144 639344 386196 639396
rect 397920 639344 397972 639396
rect 398840 639344 398892 639396
rect 400220 639276 400272 639328
rect 402336 639208 402388 639260
rect 401968 639140 402020 639192
rect 400404 639072 400456 639124
rect 402520 639004 402572 639056
rect 403900 638936 403952 638988
rect 49424 636692 49476 636744
rect 50528 636692 50580 636744
rect 403624 634788 403676 634840
rect 478696 634788 478748 634840
rect 254400 633428 254452 633480
rect 271236 633428 271288 633480
rect 523684 632000 523736 632052
rect 580172 632000 580224 632052
rect 49148 629348 49200 629400
rect 50436 629348 50488 629400
rect 254308 627920 254360 627972
rect 278044 627920 278096 627972
rect 254032 622412 254084 622464
rect 264244 622412 264296 622464
rect 48780 619012 48832 619064
rect 50344 619012 50396 619064
rect 538864 616836 538916 616888
rect 580172 616836 580224 616888
rect 254492 611328 254544 611380
rect 269764 611328 269816 611380
rect 254216 604460 254268 604512
rect 275284 604460 275336 604512
rect 398380 600244 398432 600296
rect 403624 600244 403676 600296
rect 364800 600176 364852 600228
rect 365168 600176 365220 600228
rect 300952 599836 301004 599888
rect 302194 599836 302246 599888
rect 306380 599836 306432 599888
rect 307714 599836 307766 599888
rect 382280 599836 382332 599888
rect 400588 599836 400640 599888
rect 379796 599768 379848 599820
rect 399208 599768 399260 599820
rect 378416 599700 378468 599752
rect 399300 599700 399352 599752
rect 372620 599632 372672 599684
rect 399392 599632 399444 599684
rect 365720 599564 365772 599616
rect 400496 599564 400548 599616
rect 300860 599360 300912 599412
rect 301412 599360 301464 599412
rect 357072 599360 357124 599412
rect 283012 599292 283064 599344
rect 333244 599292 333296 599344
rect 305000 599224 305052 599276
rect 305920 599224 305972 599276
rect 355600 599224 355652 599276
rect 302148 599156 302200 599208
rect 353208 599156 353260 599208
rect 359648 599156 359700 599208
rect 360016 599156 360068 599208
rect 404728 599156 404780 599208
rect 296720 599088 296772 599140
rect 298008 599088 298060 599140
rect 349896 599088 349948 599140
rect 387708 599088 387760 599140
rect 405004 599088 405056 599140
rect 353116 599020 353168 599072
rect 361580 599020 361632 599072
rect 361764 599020 361816 599072
rect 472624 599020 472676 599072
rect 254124 598952 254176 599004
rect 273904 598952 273956 599004
rect 299480 598952 299532 599004
rect 300308 598952 300360 599004
rect 361028 598952 361080 599004
rect 386604 598952 386656 599004
rect 387708 598952 387760 599004
rect 299388 598884 299440 598936
rect 359648 598884 359700 598936
rect 388260 598884 388312 598936
rect 521752 598884 521804 598936
rect 304724 598816 304776 598868
rect 361212 598816 361264 598868
rect 386420 598816 386472 598868
rect 387156 598816 387208 598868
rect 513840 598816 513892 598868
rect 298652 598748 298704 598800
rect 299388 598748 299440 598800
rect 355508 598748 355560 598800
rect 388444 598748 388496 598800
rect 478144 598748 478196 598800
rect 305828 598680 305880 598732
rect 306288 598680 306340 598732
rect 361120 598680 361172 598732
rect 304172 598612 304224 598664
rect 304632 598612 304684 598664
rect 357164 598612 357216 598664
rect 361028 598612 361080 598664
rect 381084 598612 381136 598664
rect 304908 598544 304960 598596
rect 342904 598544 342956 598596
rect 363604 598544 363656 598596
rect 371700 598544 371752 598596
rect 377220 598544 377272 598596
rect 397644 598544 397696 598596
rect 294512 598476 294564 598528
rect 300124 598476 300176 598528
rect 308312 598476 308364 598528
rect 357072 598476 357124 598528
rect 366180 598476 366232 598528
rect 397736 598476 397788 598528
rect 317328 598408 317380 598460
rect 401048 598408 401100 598460
rect 290924 598340 290976 598392
rect 404636 598340 404688 598392
rect 288992 598272 289044 598324
rect 403256 598272 403308 598324
rect 284576 598204 284628 598256
rect 403348 598204 403400 598256
rect 471244 598204 471296 598256
rect 496452 598204 496504 598256
rect 282920 598136 282972 598188
rect 283656 598136 283708 598188
rect 285588 598136 285640 598188
rect 286324 598136 286376 598188
rect 291108 598136 291160 598188
rect 291844 598136 291896 598188
rect 292580 598136 292632 598188
rect 293592 598136 293644 598188
rect 295340 598136 295392 598188
rect 295800 598136 295852 598188
rect 299204 598136 299256 598188
rect 300676 598136 300728 598188
rect 302884 598136 302936 598188
rect 311072 598136 311124 598188
rect 311992 598136 312044 598188
rect 312912 598136 312964 598188
rect 313280 598136 313332 598188
rect 314016 598136 314068 598188
rect 314660 598136 314712 598188
rect 315120 598136 315172 598188
rect 316868 598136 316920 598188
rect 324964 598136 325016 598188
rect 364432 598136 364484 598188
rect 365260 598136 365312 598188
rect 367100 598136 367152 598188
rect 368020 598136 368072 598188
rect 372804 598136 372856 598188
rect 372988 598136 373040 598188
rect 376668 598136 376720 598188
rect 377404 598136 377456 598188
rect 378324 598136 378376 598188
rect 379060 598136 379112 598188
rect 379612 598136 379664 598188
rect 380164 598136 380216 598188
rect 380992 598136 381044 598188
rect 381820 598136 381872 598188
rect 382372 598136 382424 598188
rect 382924 598136 382976 598188
rect 385040 598136 385092 598188
rect 385684 598136 385736 598188
rect 388260 598136 388312 598188
rect 388536 598136 388588 598188
rect 389272 598136 389324 598188
rect 390100 598136 390152 598188
rect 393320 598136 393372 598188
rect 393964 598136 394016 598188
rect 394700 598136 394752 598188
rect 395068 598136 395120 598188
rect 396080 598136 396132 598188
rect 396724 598136 396776 598188
rect 291200 598068 291252 598120
rect 291936 598068 291988 598120
rect 309140 598068 309192 598120
rect 310152 598068 310204 598120
rect 311900 598068 311952 598120
rect 312360 598068 312412 598120
rect 372712 598068 372764 598120
rect 373540 598068 373592 598120
rect 300768 598000 300820 598052
rect 319536 598000 319588 598052
rect 290372 597796 290424 597848
rect 294604 597796 294656 597848
rect 286876 597592 286928 597644
rect 289084 597592 289136 597644
rect 390560 597592 390612 597644
rect 391204 597592 391256 597644
rect 327724 596912 327776 596964
rect 311072 596844 311124 596896
rect 336004 596844 336056 596896
rect 342168 596844 342220 596896
rect 363972 596844 364024 596896
rect 297548 596776 297600 596828
rect 327724 596776 327776 596828
rect 329104 596776 329156 596828
rect 398196 596776 398248 596828
rect 384396 596572 384448 596624
rect 392584 596572 392636 596624
rect 302240 595552 302292 595604
rect 334624 595552 334676 595604
rect 362960 595552 363012 595604
rect 387800 595552 387852 595604
rect 333888 595484 333940 595536
rect 367376 595484 367428 595536
rect 291292 595416 291344 595468
rect 345664 595416 345716 595468
rect 347780 595416 347832 595468
rect 510712 595416 510764 595468
rect 49516 594804 49568 594856
rect 51816 594804 51868 594856
rect 288072 594192 288124 594244
rect 331956 594192 332008 594244
rect 324228 594124 324280 594176
rect 375380 594124 375432 594176
rect 381544 594124 381596 594176
rect 386420 594124 386472 594176
rect 311164 594056 311216 594108
rect 327816 594056 327868 594108
rect 331220 594056 331272 594108
rect 499580 594056 499632 594108
rect 254768 593376 254820 593428
rect 271144 593376 271196 593428
rect 266360 592628 266412 592680
rect 498200 592628 498252 592680
rect 312084 591948 312136 592000
rect 316684 591948 316736 592000
rect 325516 591336 325568 591388
rect 364708 591336 364760 591388
rect 371884 591336 371936 591388
rect 392032 591336 392084 591388
rect 293960 591268 294012 591320
rect 386788 591268 386840 591320
rect 485872 590656 485924 590708
rect 579804 590656 579856 590708
rect 49608 590588 49660 590640
rect 51724 590588 51776 590640
rect 306748 589976 306800 590028
rect 333244 589976 333296 590028
rect 336648 589976 336700 590028
rect 369032 589976 369084 590028
rect 292948 589908 293000 589960
rect 349896 589908 349948 589960
rect 361120 589908 361172 589960
rect 391940 589908 391992 589960
rect 385684 589228 385736 589280
rect 390652 589228 390704 589280
rect 311992 588616 312044 588668
rect 338856 588616 338908 588668
rect 343548 588616 343600 588668
rect 371792 588616 371844 588668
rect 288440 588548 288492 588600
rect 347044 588548 347096 588600
rect 254492 587936 254544 587988
rect 260104 587936 260156 587988
rect 329288 587120 329340 587172
rect 372896 587120 372948 587172
rect 322480 585760 322532 585812
rect 506480 585760 506532 585812
rect 340144 584536 340196 584588
rect 396172 584536 396224 584588
rect 307760 584468 307812 584520
rect 368572 584468 368624 584520
rect 287152 584400 287204 584452
rect 353116 584400 353168 584452
rect 285680 582972 285732 583024
rect 347136 582972 347188 583024
rect 385776 582360 385828 582412
rect 389272 582360 389324 582412
rect 253940 581272 253992 581324
rect 255964 581272 256016 581324
rect 310520 580252 310572 580304
rect 374276 580252 374328 580304
rect 322388 578144 322440 578196
rect 580172 578144 580224 578196
rect 300860 577464 300912 577516
rect 342904 577464 342956 577516
rect 314844 576172 314896 576224
rect 390652 576172 390704 576224
rect 286324 576104 286376 576156
rect 386604 576104 386656 576156
rect 254492 575492 254544 575544
rect 261484 575492 261536 575544
rect 323676 574744 323728 574796
rect 382464 574744 382516 574796
rect 313372 573384 313424 573436
rect 376944 573384 376996 573436
rect 292580 573316 292632 573368
rect 357164 573316 357216 573368
rect 306380 571956 306432 572008
rect 389272 571956 389324 572008
rect 283012 570664 283064 570716
rect 350080 570664 350132 570716
rect 304724 570596 304776 570648
rect 394884 570596 394936 570648
rect 253940 569984 253992 570036
rect 256056 569984 256108 570036
rect 314752 569236 314804 569288
rect 337476 569236 337528 569288
rect 253388 569168 253440 569220
rect 512092 569168 512144 569220
rect 388628 568556 388680 568608
rect 393412 568556 393464 568608
rect 355876 567808 355928 567860
rect 367100 567808 367152 567860
rect 358176 566516 358228 566568
rect 394792 566516 394844 566568
rect 305000 566448 305052 566500
rect 365904 566448 365956 566500
rect 385132 565496 385184 565548
rect 391940 565496 391992 565548
rect 296720 565156 296772 565208
rect 367376 565156 367428 565208
rect 253296 565088 253348 565140
rect 381084 565088 381136 565140
rect 300124 563728 300176 563780
rect 367192 563728 367244 563780
rect 254584 563660 254636 563712
rect 320180 563660 320232 563712
rect 359096 563660 359148 563712
rect 380992 563660 381044 563712
rect 358084 562436 358136 562488
rect 390560 562436 390612 562488
rect 300768 562368 300820 562420
rect 363052 562368 363104 562420
rect 372804 562368 372856 562420
rect 383844 562368 383896 562420
rect 291844 562300 291896 562352
rect 375380 562300 375432 562352
rect 321100 561076 321152 561128
rect 402152 561076 402204 561128
rect 304816 561008 304868 561060
rect 399944 561008 399996 561060
rect 289084 560940 289136 560992
rect 386696 560940 386748 560992
rect 362960 559648 363012 559700
rect 374092 559648 374144 559700
rect 358268 559580 358320 559632
rect 386512 559580 386564 559632
rect 265624 559512 265676 559564
rect 483112 559512 483164 559564
rect 365812 558832 365864 558884
rect 371608 558832 371660 558884
rect 359004 558288 359056 558340
rect 381176 558288 381228 558340
rect 362592 558220 362644 558272
rect 374000 558220 374052 558272
rect 376852 558220 376904 558272
rect 538864 558220 538916 558272
rect 264336 558152 264388 558204
rect 512276 558152 512328 558204
rect 254584 557540 254636 557592
rect 265624 557540 265676 557592
rect 372712 557540 372764 557592
rect 404360 557540 404412 557592
rect 355232 556996 355284 557048
rect 372712 556996 372764 557048
rect 359372 556860 359424 556912
rect 379612 556860 379664 556912
rect 358360 556792 358412 556844
rect 396080 556792 396132 556844
rect 359280 555500 359332 555552
rect 385040 555500 385092 555552
rect 253204 555432 253256 555484
rect 512000 555432 512052 555484
rect 369860 554752 369912 554804
rect 403072 554752 403124 554804
rect 355692 554072 355744 554124
rect 369860 554072 369912 554124
rect 295524 554004 295576 554056
rect 404820 554004 404872 554056
rect 358728 553392 358780 553444
rect 361028 553392 361080 553444
rect 376852 553324 376904 553376
rect 377772 553324 377824 553376
rect 392584 553324 392636 553376
rect 394148 553324 394200 553376
rect 360108 553052 360160 553104
rect 378692 553052 378744 553104
rect 356888 552984 356940 553036
rect 376760 552984 376812 553036
rect 392860 552984 392912 553036
rect 398932 552984 398984 553036
rect 356980 552916 357032 552968
rect 396356 552916 396408 552968
rect 322296 552848 322348 552900
rect 364524 552848 364576 552900
rect 389640 552848 389692 552900
rect 400404 552848 400456 552900
rect 309232 552780 309284 552832
rect 360660 552780 360712 552832
rect 361488 552780 361540 552832
rect 374184 552780 374236 552832
rect 376116 552780 376168 552832
rect 399024 552780 399076 552832
rect 322204 552712 322256 552764
rect 380624 552712 380676 552764
rect 383752 552712 383804 552764
rect 399484 552712 399536 552764
rect 325056 552644 325108 552696
rect 397368 552644 397420 552696
rect 393504 552440 393556 552492
rect 399116 552440 399168 552492
rect 356060 552372 356112 552424
rect 371884 552372 371936 552424
rect 355784 552304 355836 552356
rect 381544 552304 381596 552356
rect 354956 552236 355008 552288
rect 385776 552372 385828 552424
rect 348424 552168 348476 552220
rect 387984 552304 388036 552356
rect 396724 552236 396776 552288
rect 398012 552236 398064 552288
rect 398656 552236 398708 552288
rect 418804 552236 418856 552288
rect 384488 552168 384540 552220
rect 385684 552168 385736 552220
rect 394792 552168 394844 552220
rect 430580 552168 430632 552220
rect 367100 552100 367152 552152
rect 414664 552100 414716 552152
rect 373540 552032 373592 552084
rect 420184 552032 420236 552084
rect 393320 551964 393372 552016
rect 400588 551964 400640 552016
rect 389180 551692 389232 551744
rect 399852 551692 399904 551744
rect 383660 551624 383712 551676
rect 400036 551624 400088 551676
rect 363236 551556 363288 551608
rect 400404 551556 400456 551608
rect 360108 551488 360160 551540
rect 444380 551488 444432 551540
rect 295340 551420 295392 551472
rect 402980 551420 403032 551472
rect 295432 551352 295484 551404
rect 404452 551352 404504 551404
rect 254400 551284 254452 551336
rect 268384 551284 268436 551336
rect 291200 551284 291252 551336
rect 403440 551284 403492 551336
rect 382280 551216 382332 551268
rect 382924 551216 382976 551268
rect 354220 551080 354272 551132
rect 388628 551080 388680 551132
rect 388996 551080 389048 551132
rect 377404 551012 377456 551064
rect 377956 551012 378008 551064
rect 403532 551012 403584 551064
rect 351460 550944 351512 550996
rect 384488 550944 384540 550996
rect 355508 550876 355560 550928
rect 397460 550876 397512 550928
rect 355600 550808 355652 550860
rect 404544 550808 404596 550860
rect 345848 550740 345900 550792
rect 364432 550740 364484 550792
rect 396080 550740 396132 550792
rect 333336 550672 333388 550724
rect 333888 550672 333940 550724
rect 404912 550672 404964 550724
rect 356980 550604 357032 550656
rect 361120 550604 361172 550656
rect 391204 550604 391256 550656
rect 475844 550604 475896 550656
rect 399760 550536 399812 550588
rect 402060 550536 402112 550588
rect 397552 550468 397604 550520
rect 400680 550468 400732 550520
rect 386604 550264 386656 550316
rect 387064 550264 387116 550316
rect 356888 550128 356940 550180
rect 362960 550128 363012 550180
rect 355140 550060 355192 550112
rect 362592 550060 362644 550112
rect 352472 549992 352524 550044
rect 377956 549992 378008 550044
rect 355048 549924 355100 549976
rect 394700 549992 394752 550044
rect 400772 549992 400824 550044
rect 322204 549856 322256 549908
rect 397644 549856 397696 549908
rect 402428 549856 402480 549908
rect 364892 549788 364944 549840
rect 371332 549788 371384 549840
rect 345756 549380 345808 549432
rect 353208 549448 353260 549500
rect 326988 549312 327040 549364
rect 355140 549312 355192 549364
rect 325056 549244 325108 549296
rect 383660 549788 383712 549840
rect 322296 548564 322348 548616
rect 356060 548564 356112 548616
rect 304908 548496 304960 548548
rect 341524 548496 341576 548548
rect 281540 547816 281592 547868
rect 357440 547816 357492 547868
rect 316684 546388 316736 546440
rect 357440 546388 357492 546440
rect 279516 545844 279568 545896
rect 313648 545844 313700 545896
rect 279608 545708 279660 545760
rect 312912 545708 312964 545760
rect 313280 545708 313332 545760
rect 349988 545708 350040 545760
rect 307668 545028 307720 545080
rect 357440 545028 357492 545080
rect 278964 543600 279016 543652
rect 297456 543600 297508 543652
rect 279240 543532 279292 543584
rect 300400 543532 300452 543584
rect 279976 543464 280028 543516
rect 301136 543464 301188 543516
rect 280068 543396 280120 543448
rect 302608 543396 302660 543448
rect 401600 543396 401652 543448
rect 404544 543396 404596 543448
rect 279424 543328 279476 543380
rect 303804 543328 303856 543380
rect 279332 543260 279384 543312
rect 305552 543260 305604 543312
rect 279148 543192 279200 543244
rect 316040 543192 316092 543244
rect 279056 543124 279108 543176
rect 315120 543124 315172 543176
rect 278136 543056 278188 543108
rect 316592 543056 316644 543108
rect 257436 542988 257488 543040
rect 314844 542988 314896 543040
rect 323676 542988 323728 543040
rect 357532 542988 357584 543040
rect 279700 542580 279752 542632
rect 294512 542580 294564 542632
rect 279608 542512 279660 542564
rect 293960 542512 294012 542564
rect 279884 542444 279936 542496
rect 295340 542444 295392 542496
rect 279516 542376 279568 542428
rect 295984 542376 296036 542428
rect 306288 541696 306340 541748
rect 340236 541696 340288 541748
rect 254676 541628 254728 541680
rect 267004 541628 267056 541680
rect 309140 541628 309192 541680
rect 354128 541628 354180 541680
rect 254584 541152 254636 541204
rect 260196 541152 260248 541204
rect 401600 540948 401652 541000
rect 437480 540948 437532 541000
rect 317420 540200 317472 540252
rect 330484 540200 330536 540252
rect 278320 539656 278372 539708
rect 283472 539656 283524 539708
rect 276664 539588 276716 539640
rect 286416 539588 286468 539640
rect 280804 539520 280856 539572
rect 284208 539520 284260 539572
rect 330484 539520 330536 539572
rect 357440 539520 357492 539572
rect 281172 539452 281224 539504
rect 284944 539452 284996 539504
rect 320180 537480 320232 537532
rect 325608 537480 325660 537532
rect 329104 537480 329156 537532
rect 340880 536800 340932 536852
rect 358360 536800 358412 536852
rect 485504 536800 485556 536852
rect 579896 536800 579948 536852
rect 349896 536732 349948 536784
rect 357440 536732 357492 536784
rect 355416 536664 355468 536716
rect 357900 536664 357952 536716
rect 401600 536188 401652 536240
rect 403348 536188 403400 536240
rect 322388 536052 322440 536104
rect 340880 536052 340932 536104
rect 477500 536052 477552 536104
rect 502892 536052 502944 536104
rect 338856 535372 338908 535424
rect 357440 535372 357492 535424
rect 350080 535304 350132 535356
rect 357532 535304 357584 535356
rect 353116 535236 353168 535288
rect 357440 535236 357492 535288
rect 322480 534692 322532 534744
rect 330484 534692 330536 534744
rect 254676 534080 254728 534132
rect 278136 534080 278188 534132
rect 322480 534080 322532 534132
rect 359740 534080 359792 534132
rect 401876 533740 401928 533792
rect 404360 533740 404412 533792
rect 358176 533468 358228 533520
rect 322848 533400 322900 533452
rect 340144 533400 340196 533452
rect 328368 533332 328420 533384
rect 357716 533332 357768 533384
rect 481548 533332 481600 533384
rect 526444 533332 526496 533384
rect 323768 532720 323820 532772
rect 350540 532720 350592 532772
rect 321652 532652 321704 532704
rect 355140 532652 355192 532704
rect 327816 532584 327868 532636
rect 357440 532584 357492 532636
rect 336004 532516 336056 532568
rect 357532 532516 357584 532568
rect 350540 532448 350592 532500
rect 351184 532448 351236 532500
rect 355232 532448 355284 532500
rect 475476 531972 475528 532024
rect 492680 531972 492732 532024
rect 494428 531972 494480 532024
rect 582380 531972 582432 532024
rect 401968 531904 402020 531956
rect 404728 531904 404780 531956
rect 434720 531904 434772 531956
rect 505560 531904 505612 531956
rect 416780 531836 416832 531888
rect 497740 531836 497792 531888
rect 438860 531768 438912 531820
rect 496452 531768 496504 531820
rect 475384 531700 475436 531752
rect 506112 531700 506164 531752
rect 507216 531700 507268 531752
rect 549904 531700 549956 531752
rect 476764 531632 476816 531684
rect 508780 531632 508832 531684
rect 463700 531564 463752 531616
rect 495440 531564 495492 531616
rect 499304 531564 499356 531616
rect 527824 531564 527876 531616
rect 448520 531496 448572 531548
rect 487436 531496 487488 531548
rect 504180 531496 504232 531548
rect 534724 531496 534776 531548
rect 476948 531428 477000 531480
rect 488080 531428 488132 531480
rect 508688 531428 508740 531480
rect 538864 531428 538916 531480
rect 473360 531360 473412 531412
rect 486792 531360 486844 531412
rect 493876 531360 493928 531412
rect 509884 531360 509936 531412
rect 476856 531292 476908 531344
rect 483572 531292 483624 531344
rect 505468 531292 505520 531344
rect 510620 531292 510672 531344
rect 401968 531224 402020 531276
rect 404452 531224 404504 531276
rect 322480 531156 322532 531208
rect 328368 531156 328420 531208
rect 485044 530544 485096 530596
rect 491944 530544 491996 530596
rect 407120 530476 407172 530528
rect 495808 530476 495860 530528
rect 475568 530408 475620 530460
rect 494520 530408 494572 530460
rect 478880 530340 478932 530392
rect 500316 530340 500368 530392
rect 357716 530272 357768 530324
rect 359464 530272 359516 530324
rect 468484 530272 468536 530324
rect 485044 530272 485096 530324
rect 472624 530204 472676 530256
rect 497096 530204 497148 530256
rect 485826 530136 485878 530188
rect 563060 530136 563112 530188
rect 409880 530068 409932 530120
rect 491622 530068 491674 530120
rect 322388 529932 322440 529984
rect 359832 530000 359884 530052
rect 402888 530000 402940 530052
rect 458180 530000 458232 530052
rect 480996 530000 481048 530052
rect 565820 530000 565872 530052
rect 400864 529932 400916 529984
rect 401876 529932 401928 529984
rect 491208 529932 491260 529984
rect 571984 529932 572036 529984
rect 322480 529864 322532 529916
rect 354220 529864 354272 529916
rect 406384 529864 406436 529916
rect 477500 529864 477552 529916
rect 337476 529796 337528 529848
rect 357440 529796 357492 529848
rect 322848 529184 322900 529236
rect 337568 529184 337620 529236
rect 509792 528844 509844 528896
rect 513380 528844 513432 528896
rect 254216 528572 254268 528624
rect 269856 528572 269908 528624
rect 402888 528572 402940 528624
rect 409144 528572 409196 528624
rect 416044 528572 416096 528624
rect 477500 528572 477552 528624
rect 513288 528572 513340 528624
rect 518164 528572 518216 528624
rect 322480 528504 322532 528556
rect 356980 528504 357032 528556
rect 401968 528300 402020 528352
rect 404636 528300 404688 528352
rect 509884 527824 509936 527876
rect 569960 527824 570012 527876
rect 321560 527212 321612 527264
rect 323676 527212 323728 527264
rect 420920 527144 420972 527196
rect 477500 527144 477552 527196
rect 322480 527076 322532 527128
rect 351460 527076 351512 527128
rect 355324 527076 355376 527128
rect 357900 527076 357952 527128
rect 331864 527008 331916 527060
rect 357440 527008 357492 527060
rect 402244 526736 402296 526788
rect 405096 526736 405148 526788
rect 401784 526396 401836 526448
rect 478880 526396 478932 526448
rect 405096 525784 405148 525836
rect 477500 525784 477552 525836
rect 322480 525716 322532 525768
rect 355048 525716 355100 525768
rect 399668 525716 399720 525768
rect 402428 525716 402480 525768
rect 422944 525716 422996 525768
rect 478696 525716 478748 525768
rect 530584 525716 530636 525768
rect 580172 525716 580224 525768
rect 475752 525580 475804 525632
rect 477960 525580 478012 525632
rect 402244 525308 402296 525360
rect 404912 525308 404964 525360
rect 322756 525036 322808 525088
rect 349896 525036 349948 525088
rect 512644 524424 512696 524476
rect 525064 524424 525116 524476
rect 333244 524356 333296 524408
rect 357440 524356 357492 524408
rect 471336 523200 471388 523252
rect 477500 523200 477552 523252
rect 254032 522996 254084 523048
rect 275376 522996 275428 523048
rect 322480 522996 322532 523048
rect 355876 522996 355928 523048
rect 456800 522996 456852 523048
rect 477500 522996 477552 523048
rect 322020 522928 322072 522980
rect 355784 522928 355836 522980
rect 357624 522928 357676 522980
rect 359648 522928 359700 522980
rect 322480 521636 322532 521688
rect 351460 521636 351512 521688
rect 402888 521636 402940 521688
rect 423680 521636 423732 521688
rect 322020 521568 322072 521620
rect 352472 521568 352524 521620
rect 352472 521024 352524 521076
rect 353300 521024 353352 521076
rect 401600 520956 401652 521008
rect 403532 520956 403584 521008
rect 322480 520276 322532 520328
rect 353116 520276 353168 520328
rect 450544 520276 450596 520328
rect 477500 520276 477552 520328
rect 353024 520208 353076 520260
rect 357440 520208 357492 520260
rect 401600 520140 401652 520192
rect 403808 520140 403860 520192
rect 322848 519528 322900 519580
rect 324228 519528 324280 519580
rect 355416 519528 355468 519580
rect 321560 519256 321612 519308
rect 323676 519256 323728 519308
rect 454684 518916 454736 518968
rect 478512 518916 478564 518968
rect 513288 518916 513340 518968
rect 531964 518916 532016 518968
rect 321836 518848 321888 518900
rect 325700 518848 325752 518900
rect 345664 518848 345716 518900
rect 357440 518848 357492 518900
rect 322480 517556 322532 517608
rect 350540 517556 350592 517608
rect 356888 517556 356940 517608
rect 466460 517556 466512 517608
rect 477592 517556 477644 517608
rect 254492 517488 254544 517540
rect 274088 517488 274140 517540
rect 326344 517488 326396 517540
rect 357532 517488 357584 517540
rect 436744 517488 436796 517540
rect 477500 517488 477552 517540
rect 321560 517420 321612 517472
rect 323768 517420 323820 517472
rect 341524 517420 341576 517472
rect 357440 517420 357492 517472
rect 477132 517420 477184 517472
rect 478512 517420 478564 517472
rect 322388 516740 322440 516792
rect 356888 516672 356940 516724
rect 322388 516332 322440 516384
rect 322940 516332 322992 516384
rect 325056 516332 325108 516384
rect 513196 516196 513248 516248
rect 526444 516196 526496 516248
rect 402612 516128 402664 516180
rect 405924 516128 405976 516180
rect 513288 516128 513340 516180
rect 536104 516128 536156 516180
rect 321836 516060 321888 516112
rect 342260 516060 342312 516112
rect 401600 516060 401652 516112
rect 403440 516060 403492 516112
rect 513196 516060 513248 516112
rect 520924 516060 520976 516112
rect 322848 515380 322900 515432
rect 324228 515380 324280 515432
rect 329288 515380 329340 515432
rect 342260 515380 342312 515432
rect 343548 515380 343600 515432
rect 353024 515380 353076 515432
rect 358084 514836 358136 514888
rect 359556 514836 359608 514888
rect 331956 514700 332008 514752
rect 357440 514700 357492 514752
rect 322112 514020 322164 514072
rect 332048 514020 332100 514072
rect 460204 513408 460256 513460
rect 477592 513408 477644 513460
rect 322480 513340 322532 513392
rect 355324 513340 355376 513392
rect 441620 513340 441672 513392
rect 477500 513340 477552 513392
rect 320364 513272 320416 513324
rect 355692 513272 355744 513324
rect 358268 513272 358320 513324
rect 359464 513272 359516 513324
rect 412640 513272 412692 513324
rect 477592 513272 477644 513324
rect 329196 513204 329248 513256
rect 357440 513204 357492 513256
rect 402520 513204 402572 513256
rect 405740 513204 405792 513256
rect 322112 512592 322164 512644
rect 357164 512592 357216 512644
rect 340236 511912 340288 511964
rect 357440 511912 357492 511964
rect 321560 511232 321612 511284
rect 336648 511232 336700 511284
rect 356980 511232 357032 511284
rect 320364 510824 320416 510876
rect 320640 510824 320692 510876
rect 327908 510824 327960 510876
rect 254400 510620 254452 510672
rect 271328 510620 271380 510672
rect 402888 510620 402940 510672
rect 451280 510620 451332 510672
rect 462964 510620 463016 510672
rect 477592 510620 477644 510672
rect 513288 510620 513340 510672
rect 544384 510620 544436 510672
rect 320088 510552 320140 510604
rect 355600 510552 355652 510604
rect 462320 510552 462372 510604
rect 477500 510552 477552 510604
rect 320456 510484 320508 510536
rect 333336 510484 333388 510536
rect 337568 510484 337620 510536
rect 357440 510484 357492 510536
rect 324228 509872 324280 509924
rect 350080 509872 350132 509924
rect 402888 509328 402940 509380
rect 404912 509328 404964 509380
rect 445024 509328 445076 509380
rect 422944 509260 422996 509312
rect 477500 509260 477552 509312
rect 513288 509260 513340 509312
rect 522304 509260 522356 509312
rect 320180 509192 320232 509244
rect 353208 509192 353260 509244
rect 342904 509124 342956 509176
rect 357532 509124 357584 509176
rect 347044 509056 347096 509108
rect 357440 509056 357492 509108
rect 478788 508444 478840 508496
rect 479524 508444 479576 508496
rect 319076 508240 319128 508292
rect 319352 508240 319404 508292
rect 50804 507832 50856 507884
rect 51172 507832 51224 507884
rect 319076 507832 319128 507884
rect 357164 507832 357216 507884
rect 358728 507832 358780 507884
rect 359740 507832 359792 507884
rect 320364 507764 320416 507816
rect 355508 507764 355560 507816
rect 334624 507696 334676 507748
rect 357440 507696 357492 507748
rect 320088 507628 320140 507680
rect 345848 507628 345900 507680
rect 318984 506472 319036 506524
rect 320088 506472 320140 506524
rect 320180 506404 320232 506456
rect 345756 506404 345808 506456
rect 347136 506404 347188 506456
rect 357440 506404 357492 506456
rect 402244 506404 402296 506456
rect 404820 506404 404872 506456
rect 349988 506336 350040 506388
rect 357532 506336 357584 506388
rect 319352 505724 319404 505776
rect 325516 505724 325568 505776
rect 356612 505724 356664 505776
rect 318892 505520 318944 505572
rect 319352 505520 319404 505572
rect 472716 505520 472768 505572
rect 477500 505520 477552 505572
rect 254308 505112 254360 505164
rect 275468 505112 275520 505164
rect 320180 505112 320232 505164
rect 320732 505112 320784 505164
rect 340880 505112 340932 505164
rect 342168 505112 342220 505164
rect 359740 505112 359792 505164
rect 405004 505112 405056 505164
rect 477500 505112 477552 505164
rect 327724 505044 327776 505096
rect 357440 505044 357492 505096
rect 320088 504976 320140 505028
rect 340880 504976 340932 505028
rect 322388 504160 322440 504212
rect 326344 504160 326396 504212
rect 436836 503752 436888 503804
rect 477592 503752 477644 503804
rect 400864 503684 400916 503736
rect 477500 503684 477552 503736
rect 513288 503684 513340 503736
rect 530584 503684 530636 503736
rect 320180 503616 320232 503668
rect 325608 503616 325660 503668
rect 357440 503616 357492 503668
rect 401692 503616 401744 503668
rect 405832 503616 405884 503668
rect 322388 503548 322440 503600
rect 348424 503548 348476 503600
rect 478512 502596 478564 502648
rect 478788 502596 478840 502648
rect 322388 502324 322440 502376
rect 355508 502324 355560 502376
rect 440884 502324 440936 502376
rect 477500 502324 477552 502376
rect 513288 502324 513340 502376
rect 545764 502324 545816 502376
rect 337384 502256 337436 502308
rect 357440 502256 357492 502308
rect 402244 500964 402296 501016
rect 477500 500964 477552 501016
rect 352564 500896 352616 500948
rect 399484 500896 399536 500948
rect 478604 500896 478656 500948
rect 510712 500896 510764 500948
rect 353116 500828 353168 500880
rect 402060 500828 402112 500880
rect 358360 500760 358412 500812
rect 359372 500760 359424 500812
rect 510712 500760 510764 500812
rect 510988 500760 511040 500812
rect 510988 500624 511040 500676
rect 511264 500624 511316 500676
rect 296628 500352 296680 500404
rect 321744 500352 321796 500404
rect 295248 500284 295300 500336
rect 321652 500284 321704 500336
rect 292764 500216 292816 500268
rect 320640 500216 320692 500268
rect 322204 500216 322256 500268
rect 360844 499944 360896 499996
rect 254216 499876 254268 499928
rect 257436 499876 257488 499928
rect 401876 499536 401928 499588
rect 433340 499536 433392 499588
rect 468576 499536 468628 499588
rect 477500 499536 477552 499588
rect 355968 499468 356020 499520
rect 364524 499468 364576 499520
rect 394148 499468 394200 499520
rect 403716 499468 403768 499520
rect 478788 499468 478840 499520
rect 482376 499468 482428 499520
rect 373540 499400 373592 499452
rect 471244 499400 471296 499452
rect 487804 499400 487856 499452
rect 525156 499400 525208 499452
rect 322296 499332 322348 499384
rect 400772 499332 400824 499384
rect 477040 499332 477092 499384
rect 499304 499332 499356 499384
rect 353024 499264 353076 499316
rect 398012 499264 398064 499316
rect 492312 499264 492364 499316
rect 511356 499264 511408 499316
rect 359832 499196 359884 499248
rect 401692 499196 401744 499248
rect 359740 499128 359792 499180
rect 401600 499128 401652 499180
rect 359924 499060 359976 499112
rect 401968 499060 402020 499112
rect 357072 498992 357124 499044
rect 397368 498992 397420 499044
rect 356612 498924 356664 498976
rect 381912 498924 381964 498976
rect 323676 498856 323728 498908
rect 353392 498856 353444 498908
rect 367744 498856 367796 498908
rect 254584 498788 254636 498840
rect 282184 498788 282236 498840
rect 322480 498788 322532 498840
rect 362960 498788 363012 498840
rect 508504 498788 508556 498840
rect 512000 498788 512052 498840
rect 356980 498720 357032 498772
rect 389640 498720 389692 498772
rect 479248 498720 479300 498772
rect 481640 498720 481692 498772
rect 375472 498652 375524 498704
rect 580356 498652 580408 498704
rect 324964 498584 325016 498636
rect 378048 498584 378100 498636
rect 352564 498176 352616 498228
rect 353024 498176 353076 498228
rect 478420 498176 478472 498228
rect 480904 498176 480956 498228
rect 352840 498108 352892 498160
rect 355324 498108 355376 498160
rect 355416 498108 355468 498160
rect 361304 498108 361356 498160
rect 399300 498108 399352 498160
rect 403900 498108 403952 498160
rect 475660 498108 475712 498160
rect 484492 498108 484544 498160
rect 491024 498108 491076 498160
rect 521660 498108 521712 498160
rect 357348 498040 357400 498092
rect 370964 498040 371016 498092
rect 396724 498040 396776 498092
rect 405188 498040 405240 498092
rect 474004 498040 474056 498092
rect 503168 498040 503220 498092
rect 357256 497972 357308 498024
rect 367100 497972 367152 498024
rect 388352 497972 388404 498024
rect 405280 497972 405332 498024
rect 475844 497972 475896 498024
rect 502524 497972 502576 498024
rect 294604 497904 294656 497956
rect 316040 497904 316092 497956
rect 349804 497904 349856 497956
rect 379336 497904 379388 497956
rect 477224 497904 477276 497956
rect 496728 497904 496780 497956
rect 291936 497836 291988 497888
rect 315120 497836 315172 497888
rect 352748 497836 352800 497888
rect 379980 497836 380032 497888
rect 494796 497836 494848 497888
rect 510252 497836 510304 497888
rect 290464 497768 290516 497820
rect 327724 497768 327776 497820
rect 352932 497768 352984 497820
rect 366456 497768 366508 497820
rect 470600 497768 470652 497820
rect 485136 497768 485188 497820
rect 258724 497700 258776 497752
rect 301872 497700 301924 497752
rect 355324 497700 355376 497752
rect 363236 497700 363288 497752
rect 260288 497632 260340 497684
rect 316592 497632 316644 497684
rect 351368 497632 351420 497684
rect 394792 497632 394844 497684
rect 427820 497632 427872 497684
rect 493508 497632 493560 497684
rect 257620 497564 257672 497616
rect 317420 497564 317472 497616
rect 352656 497564 352708 497616
rect 372252 497564 372304 497616
rect 459560 497564 459612 497616
rect 505744 497564 505796 497616
rect 254676 497496 254728 497548
rect 314660 497496 314712 497548
rect 414020 497496 414072 497548
rect 492864 497496 492916 497548
rect 296536 497428 296588 497480
rect 487068 497428 487120 497480
rect 493416 497428 493468 497480
rect 507032 497428 507084 497480
rect 359372 497360 359424 497412
rect 481916 497360 481968 497412
rect 354128 497292 354180 497344
rect 383844 497292 383896 497344
rect 496176 496952 496228 497004
rect 501880 496952 501932 497004
rect 494704 496884 494756 496936
rect 498016 496884 498068 496936
rect 502340 496884 502392 496936
rect 509700 496884 509752 496936
rect 284576 496816 284628 496868
rect 286324 496816 286376 496868
rect 299848 496816 299900 496868
rect 305552 496816 305604 496868
rect 381544 496816 381596 496868
rect 384488 496816 384540 496868
rect 485044 496816 485096 496868
rect 488356 496816 488408 496868
rect 493324 496816 493376 496868
rect 494152 496816 494204 496868
rect 496084 496816 496136 496868
rect 498660 496816 498712 496868
rect 502984 496816 503036 496868
rect 503812 496816 503864 496868
rect 358176 496748 358228 496800
rect 366364 496748 366416 496800
rect 478236 496748 478288 496800
rect 482284 496748 482336 496800
rect 294144 496680 294196 496732
rect 295984 496680 296036 496732
rect 479156 496204 479208 496256
rect 488632 496204 488684 496256
rect 278780 496136 278832 496188
rect 320548 496136 320600 496188
rect 264980 496068 265032 496120
rect 320732 496068 320784 496120
rect 367100 496068 367152 496120
rect 479708 496136 479760 496188
rect 495532 496136 495584 496188
rect 552664 496136 552716 496188
rect 479340 496068 479392 496120
rect 547880 496068 547932 496120
rect 49240 495456 49292 495508
rect 50344 495456 50396 495508
rect 478328 495388 478380 495440
rect 480996 495388 481048 495440
rect 445760 494844 445812 494896
rect 512920 494844 512972 494896
rect 398840 494776 398892 494828
rect 511172 494776 511224 494828
rect 285680 494708 285732 494760
rect 320456 494708 320508 494760
rect 369124 494708 369176 494760
rect 483204 494708 483256 494760
rect 287060 494640 287112 494692
rect 287888 494640 287940 494692
rect 288440 494640 288492 494692
rect 289360 494640 289412 494692
rect 299480 494640 299532 494692
rect 300400 494640 300452 494692
rect 307760 494640 307812 494692
rect 308496 494640 308548 494692
rect 311900 494300 311952 494352
rect 312912 494300 312964 494352
rect 254584 494028 254636 494080
rect 261576 494028 261628 494080
rect 358268 493960 358320 494012
rect 362224 493960 362276 494012
rect 481088 493960 481140 494012
rect 483848 493960 483900 494012
rect 296720 493416 296772 493468
rect 297456 493416 297508 493468
rect 402980 493348 403032 493400
rect 512644 493348 512696 493400
rect 389180 493280 389232 493332
rect 510436 493280 510488 493332
rect 298836 492600 298888 492652
rect 302332 492600 302384 492652
rect 285864 491920 285916 491972
rect 292028 491920 292080 491972
rect 392216 491920 392268 491972
rect 412640 491920 412692 491972
rect 358912 489132 358964 489184
rect 580448 489132 580500 489184
rect 254676 488520 254728 488572
rect 279424 488520 279476 488572
rect 276020 487772 276072 487824
rect 320364 487772 320416 487824
rect 479064 486412 479116 486464
rect 580356 486412 580408 486464
rect 49424 485800 49476 485852
rect 51724 485800 51776 485852
rect 482376 485732 482428 485784
rect 580172 485732 580224 485784
rect 364340 482264 364392 482316
rect 497372 482264 497424 482316
rect 254400 481652 254452 481704
rect 268476 481652 268528 481704
rect 49332 481584 49384 481636
rect 50436 481584 50488 481636
rect 310612 480904 310664 480956
rect 350264 480904 350316 480956
rect 382280 480904 382332 480956
rect 506388 480904 506440 480956
rect 374000 479476 374052 479528
rect 471336 479476 471388 479528
rect 385040 478116 385092 478168
rect 460204 478116 460256 478168
rect 391940 476756 391992 476808
rect 480628 476756 480680 476808
rect 254216 476076 254268 476128
rect 265716 476076 265768 476128
rect 46388 473288 46440 473340
rect 48964 473288 49016 473340
rect 338764 471928 338816 471980
rect 580172 471928 580224 471980
rect 254492 470568 254544 470620
rect 264336 470568 264388 470620
rect 45468 467780 45520 467832
rect 48780 467780 48832 467832
rect 49056 467780 49108 467832
rect 254676 465060 254728 465112
rect 289084 465060 289136 465112
rect 47860 462272 47912 462324
rect 50804 462272 50856 462324
rect 297640 460164 297692 460216
rect 313372 460164 313424 460216
rect 254308 458192 254360 458244
rect 269948 458192 270000 458244
rect 46480 456356 46532 456408
rect 49792 456356 49844 456408
rect 299572 453976 299624 454028
rect 300952 453976 301004 454028
rect 254676 452616 254728 452668
rect 284944 452616 284996 452668
rect 50620 450712 50672 450764
rect 51264 450712 51316 450764
rect 254676 447108 254728 447160
rect 278228 447108 278280 447160
rect 46572 445680 46624 445732
rect 48320 445680 48372 445732
rect 254400 441736 254452 441788
rect 257528 441736 257580 441788
rect 46664 438812 46716 438864
rect 48320 438812 48372 438864
rect 254676 434732 254728 434784
rect 291844 434732 291896 434784
rect 46756 433236 46808 433288
rect 49148 433236 49200 433288
rect 518164 431876 518216 431928
rect 579620 431876 579672 431928
rect 254216 429156 254268 429208
rect 351460 429156 351512 429208
rect 46848 427728 46900 427780
rect 49424 427728 49476 427780
rect 254676 423648 254728 423700
rect 323676 423648 323728 423700
rect 323584 419432 323636 419484
rect 580172 419432 580224 419484
rect 254400 418140 254452 418192
rect 287704 418140 287756 418192
rect 3148 409844 3200 409896
rect 50528 409844 50580 409896
rect 254308 405696 254360 405748
rect 350816 405696 350868 405748
rect 366364 405628 366416 405680
rect 580172 405628 580224 405680
rect 254492 400188 254544 400240
rect 350632 400188 350684 400240
rect 254492 394952 254544 395004
rect 260380 394952 260432 395004
rect 46848 391960 46900 392012
rect 48320 391960 48372 392012
rect 254492 389172 254544 389224
rect 313924 389172 313976 389224
rect 46756 385024 46808 385076
rect 48320 385024 48372 385076
rect 254216 382236 254268 382288
rect 289176 382236 289228 382288
rect 46664 379516 46716 379568
rect 49424 379516 49476 379568
rect 254124 376728 254176 376780
rect 350908 376728 350960 376780
rect 254400 371220 254452 371272
rect 301504 371220 301556 371272
rect 254492 365712 254544 365764
rect 287796 365712 287848 365764
rect 320824 365644 320876 365696
rect 580172 365644 580224 365696
rect 299664 362176 299716 362228
rect 314660 362176 314712 362228
rect 253940 358844 253992 358896
rect 256148 358844 256200 358896
rect 3148 357416 3200 357468
rect 50620 357416 50672 357468
rect 307852 355308 307904 355360
rect 349804 355308 349856 355360
rect 288532 353948 288584 354000
rect 352656 353948 352708 354000
rect 482560 353948 482612 354000
rect 552020 353948 552072 354000
rect 254492 353268 254544 353320
rect 289268 353268 289320 353320
rect 362224 353200 362276 353252
rect 580172 353200 580224 353252
rect 498200 352588 498252 352640
rect 510068 352588 510120 352640
rect 287152 352520 287204 352572
rect 350172 352520 350224 352572
rect 431960 352520 432012 352572
rect 512552 352520 512604 352572
rect 289820 351160 289872 351212
rect 319168 351160 319220 351212
rect 258080 349800 258132 349852
rect 511080 349800 511132 349852
rect 299020 348372 299072 348424
rect 307760 348372 307812 348424
rect 254768 347760 254820 347812
rect 346400 347760 346452 347812
rect 288440 347012 288492 347064
rect 352104 347012 352156 347064
rect 282920 345652 282972 345704
rect 319076 345652 319128 345704
rect 3332 345040 3384 345092
rect 50252 345040 50304 345092
rect 297824 344360 297876 344412
rect 311992 344360 312044 344412
rect 271880 344292 271932 344344
rect 318984 344292 319036 344344
rect 283104 342864 283156 342916
rect 349896 342864 349948 342916
rect 254676 342252 254728 342304
rect 296168 342252 296220 342304
rect 296812 341640 296864 341692
rect 311992 341640 312044 341692
rect 303804 341572 303856 341624
rect 320272 341572 320324 341624
rect 285772 341504 285824 341556
rect 352472 341504 352524 341556
rect 478972 341504 479024 341556
rect 580356 341504 580408 341556
rect 296720 340144 296772 340196
rect 349712 340144 349764 340196
rect 267740 338784 267792 338836
rect 318892 338784 318944 338836
rect 289912 338716 289964 338768
rect 352288 338716 352340 338768
rect 299480 337492 299532 337544
rect 319352 337492 319404 337544
rect 260840 337356 260892 337408
rect 319260 337356 319312 337408
rect 254768 335996 254820 336048
rect 350724 335996 350776 336048
rect 313924 335384 313976 335436
rect 318064 335384 318116 335436
rect 254676 335316 254728 335368
rect 332232 335316 332284 335368
rect 298560 334704 298612 334756
rect 311900 334704 311952 334756
rect 310520 334636 310572 334688
rect 352012 334636 352064 334688
rect 291292 334568 291344 334620
rect 351092 334568 351144 334620
rect 306472 333344 306524 333396
rect 351000 333344 351052 333396
rect 286324 333276 286376 333328
rect 352380 333276 352432 333328
rect 298008 333208 298060 333260
rect 320180 333208 320232 333260
rect 301504 333140 301556 333192
rect 306472 333140 306524 333192
rect 285128 332188 285180 332240
rect 323216 332188 323268 332240
rect 296444 332120 296496 332172
rect 305092 332120 305144 332172
rect 349712 332120 349764 332172
rect 349988 332120 350040 332172
rect 295156 332052 295208 332104
rect 306380 332052 306432 332104
rect 296352 331984 296404 332036
rect 309140 331984 309192 332036
rect 294972 331916 295024 331968
rect 309232 331916 309284 331968
rect 295064 331848 295116 331900
rect 302424 331848 302476 331900
rect 303620 331848 303672 331900
rect 350356 331848 350408 331900
rect 323676 331780 323728 331832
rect 325148 331780 325200 331832
rect 293868 331712 293920 331764
rect 309048 331712 309100 331764
rect 298744 331644 298796 331696
rect 343824 331644 343876 331696
rect 296260 331576 296312 331628
rect 313556 331576 313608 331628
rect 292120 331508 292172 331560
rect 321928 331508 321980 331560
rect 327724 331508 327776 331560
rect 333520 331508 333572 331560
rect 338028 331508 338080 331560
rect 353576 331508 353628 331560
rect 298836 331440 298888 331492
rect 329012 331440 329064 331492
rect 339316 331440 339368 331492
rect 352196 331440 352248 331492
rect 293776 331372 293828 331424
rect 330944 331372 330996 331424
rect 336096 331372 336148 331424
rect 354680 331372 354732 331424
rect 298928 331304 298980 331356
rect 307760 331304 307812 331356
rect 327724 331304 327776 331356
rect 353668 331304 353720 331356
rect 293684 331236 293736 331288
rect 301964 331236 302016 331288
rect 345112 331236 345164 331288
rect 354772 331236 354824 331288
rect 284300 330488 284352 330540
rect 286324 330488 286376 330540
rect 299204 330080 299256 330132
rect 326436 330080 326488 330132
rect 299296 330012 299348 330064
rect 334532 330012 334584 330064
rect 299112 329944 299164 329996
rect 340236 329944 340288 329996
rect 254216 329876 254268 329928
rect 285036 329876 285088 329928
rect 299388 329876 299440 329928
rect 347412 329876 347464 329928
rect 254676 329808 254728 329860
rect 350080 329808 350132 329860
rect 254492 325592 254544 325644
rect 292120 325592 292172 325644
rect 349804 325048 349856 325100
rect 349896 325048 349948 325100
rect 349804 324844 349856 324896
rect 349896 324844 349948 324896
rect 281540 324232 281592 324284
rect 297732 324232 297784 324284
rect 254308 320084 254360 320136
rect 285128 320084 285180 320136
rect 287796 318724 287848 318776
rect 297732 318724 297784 318776
rect 285036 317364 285088 317416
rect 297732 317364 297784 317416
rect 297272 316004 297324 316056
rect 297732 316004 297784 316056
rect 351368 314644 351420 314696
rect 351920 314644 351972 314696
rect 292856 313216 292908 313268
rect 297916 313216 297968 313268
rect 354036 313216 354088 313268
rect 580172 313216 580224 313268
rect 260380 307708 260432 307760
rect 298008 307708 298060 307760
rect 254216 306348 254268 306400
rect 293316 306348 293368 306400
rect 256148 306280 256200 306332
rect 298008 306280 298060 306332
rect 349988 303628 350040 303680
rect 351920 303628 351972 303680
rect 293960 303492 294012 303544
rect 298008 303492 298060 303544
rect 292580 303152 292632 303204
rect 294696 303152 294748 303204
rect 254676 300840 254728 300892
rect 294788 300840 294840 300892
rect 383200 299412 383252 299464
rect 579620 299412 579672 299464
rect 254676 295332 254728 295384
rect 285036 295332 285088 295384
rect 297824 295128 297876 295180
rect 299756 295128 299808 295180
rect 286324 292476 286376 292528
rect 298008 292476 298060 292528
rect 295432 289620 295484 289672
rect 298008 289620 298060 289672
rect 292028 288328 292080 288380
rect 298008 288328 298060 288380
rect 297824 287376 297876 287428
rect 297824 287036 297876 287088
rect 297824 285880 297876 285932
rect 297824 285676 297876 285728
rect 289176 285608 289228 285660
rect 297916 285608 297968 285660
rect 254308 282888 254360 282940
rect 264428 282888 264480 282940
rect 3516 282004 3568 282056
rect 295432 282004 295484 282056
rect 50620 281936 50672 281988
rect 296076 281936 296128 281988
rect 46756 281868 46808 281920
rect 279884 281868 279936 281920
rect 48780 281800 48832 281852
rect 52920 281800 52972 281852
rect 3424 281460 3476 281512
rect 500592 281460 500644 281512
rect 50528 281392 50580 281444
rect 512460 281392 512512 281444
rect 49148 281324 49200 281376
rect 281172 281324 281224 281376
rect 285036 281324 285088 281376
rect 352012 281324 352064 281376
rect 48964 281256 49016 281308
rect 51908 281256 51960 281308
rect 49056 281120 49108 281172
rect 54484 281256 54536 281308
rect 55864 281256 55916 281308
rect 279792 281256 279844 281308
rect 52092 281188 52144 281240
rect 280988 281188 281040 281240
rect 48688 281052 48740 281104
rect 280804 281120 280856 281172
rect 52920 281052 52972 281104
rect 278320 281052 278372 281104
rect 49240 280984 49292 281036
rect 48044 280916 48096 280968
rect 55864 280916 55916 280968
rect 276664 280984 276716 281036
rect 254032 280916 254084 280968
rect 351460 280916 351512 280968
rect 51908 280780 51960 280832
rect 53104 280780 53156 280832
rect 297732 280576 297784 280628
rect 300124 280576 300176 280628
rect 347320 280576 347372 280628
rect 350080 280576 350132 280628
rect 50252 280100 50304 280152
rect 478144 280100 478196 280152
rect 3608 280032 3660 280084
rect 405096 280032 405148 280084
rect 46664 279964 46716 280016
rect 279700 279964 279752 280016
rect 299848 279964 299900 280016
rect 305000 279964 305052 280016
rect 46848 279896 46900 279948
rect 279516 279896 279568 279948
rect 298928 279896 298980 279948
rect 303804 279896 303856 279948
rect 48228 279828 48280 279880
rect 279608 279828 279660 279880
rect 296260 279488 296312 279540
rect 310520 279488 310572 279540
rect 59544 279420 59596 279472
rect 297364 279420 297416 279472
rect 321652 279420 321704 279472
rect 352196 279420 352248 279472
rect 289268 279012 289320 279064
rect 315488 279012 315540 279064
rect 287704 278944 287756 278996
rect 321284 278944 321336 278996
rect 296168 278876 296220 278928
rect 330944 278876 330996 278928
rect 294788 278808 294840 278860
rect 342536 278808 342588 278860
rect 293316 278740 293368 278792
rect 349620 278740 349672 278792
rect 295064 278672 295116 278724
rect 345756 278672 345808 278724
rect 296352 278604 296404 278656
rect 296444 278536 296496 278588
rect 295340 278468 295392 278520
rect 335452 278468 335504 278520
rect 294972 278400 295024 278452
rect 322572 278400 322624 278452
rect 337384 278604 337436 278656
rect 341248 278604 341300 278656
rect 339960 278468 340012 278520
rect 338028 278400 338080 278452
rect 294696 278332 294748 278384
rect 319996 278332 320048 278384
rect 295156 278264 295208 278316
rect 318064 278264 318116 278316
rect 287060 278196 287112 278248
rect 295984 278128 296036 278180
rect 300032 278196 300084 278248
rect 305644 278196 305696 278248
rect 303896 278060 303948 278112
rect 334164 278060 334216 278112
rect 338212 278060 338264 278112
rect 341524 278060 341576 278112
rect 351920 278060 351972 278112
rect 298652 277992 298704 278044
rect 303712 277992 303764 278044
rect 317420 277992 317472 278044
rect 343824 277992 343876 278044
rect 301320 277924 301372 277976
rect 308404 277924 308456 277976
rect 313280 277924 313332 277976
rect 316776 277924 316828 277976
rect 323124 277924 323176 277976
rect 323860 277516 323912 277568
rect 326344 277516 326396 277568
rect 324320 277380 324372 277432
rect 327080 277380 327132 277432
rect 297456 276700 297508 276752
rect 309140 276700 309192 276752
rect 314752 276700 314804 276752
rect 350908 276700 350960 276752
rect 8944 276632 8996 276684
rect 485780 276632 485832 276684
rect 297916 276020 297968 276072
rect 298836 276020 298888 276072
rect 297180 275340 297232 275392
rect 311164 275340 311216 275392
rect 299572 275272 299624 275324
rect 318800 275272 318852 275324
rect 297548 273912 297600 273964
rect 335360 273912 335412 273964
rect 297640 273232 297692 273284
rect 298744 273232 298796 273284
rect 479524 273164 479576 273216
rect 579896 273164 579948 273216
rect 299664 271804 299716 271856
rect 305000 271804 305052 271856
rect 13820 268404 13872 268456
rect 485044 268404 485096 268456
rect 3424 268336 3476 268388
rect 510988 268336 511040 268388
rect 301504 264188 301556 264240
rect 350724 264188 350776 264240
rect 58992 262828 59044 262880
rect 352380 262828 352432 262880
rect 58900 261468 58952 261520
rect 352748 261468 352800 261520
rect 59268 260108 59320 260160
rect 347872 260108 347924 260160
rect 356796 259360 356848 259412
rect 579804 259360 579856 259412
rect 52460 250452 52512 250504
rect 468576 250452 468628 250504
rect 359648 245556 359700 245608
rect 580172 245556 580224 245608
rect 3424 241408 3476 241460
rect 510896 241408 510948 241460
rect 9680 239368 9732 239420
rect 400864 239368 400916 239420
rect 59084 236648 59136 236700
rect 352104 236648 352156 236700
rect 57060 233928 57112 233980
rect 260288 233928 260340 233980
rect 14464 233860 14516 233912
rect 490288 233860 490340 233912
rect 486424 233180 486476 233232
rect 580172 233180 580224 233232
rect 59728 232500 59780 232552
rect 311900 232500 311952 232552
rect 59636 229712 59688 229764
rect 324412 229712 324464 229764
rect 325700 229712 325752 229764
rect 349804 229712 349856 229764
rect 57428 228352 57480 228404
rect 258724 228352 258776 228404
rect 59176 227060 59228 227112
rect 283196 227060 283248 227112
rect 308864 227060 308916 227112
rect 332600 227060 332652 227112
rect 57704 226992 57756 227044
rect 293408 226992 293460 227044
rect 318984 226992 319036 227044
rect 349712 226992 349764 227044
rect 302792 225768 302844 225820
rect 381544 225768 381596 225820
rect 58808 225700 58860 225752
rect 310612 225700 310664 225752
rect 42800 225632 42852 225684
rect 512368 225632 512420 225684
rect 3516 225564 3568 225616
rect 476948 225564 477000 225616
rect 3424 224272 3476 224324
rect 436836 224272 436888 224324
rect 3700 224204 3752 224256
rect 509884 224204 509936 224256
rect 305644 223524 305696 223576
rect 307852 223524 307904 223576
rect 311164 223524 311216 223576
rect 312912 223524 312964 223576
rect 326344 223524 326396 223576
rect 333152 223524 333204 223576
rect 300124 223456 300176 223508
rect 306840 223456 306892 223508
rect 335176 223252 335228 223304
rect 341524 223252 341576 223304
rect 302240 223184 302292 223236
rect 314936 223184 314988 223236
rect 337200 223184 337252 223236
rect 349988 223184 350040 223236
rect 309232 223116 309284 223168
rect 323032 223116 323084 223168
rect 329104 223116 329156 223168
rect 354680 223116 354732 223168
rect 299756 223048 299808 223100
rect 321008 223048 321060 223100
rect 328092 223048 328144 223100
rect 353576 223048 353628 223100
rect 293868 222980 293920 223032
rect 331128 222980 331180 223032
rect 334164 222980 334216 223032
rect 354772 222980 354824 223032
rect 57796 222912 57848 222964
rect 253572 222912 253624 222964
rect 293776 222912 293828 222964
rect 311900 222912 311952 222964
rect 316960 222912 317012 222964
rect 351368 222912 351420 222964
rect 57336 222844 57388 222896
rect 254584 222844 254636 222896
rect 293684 222844 293736 222896
rect 330116 222844 330168 222896
rect 332140 222844 332192 222896
rect 353668 222844 353720 222896
rect 222844 222232 222896 222284
rect 301504 222232 301556 222284
rect 224408 222164 224460 222216
rect 339224 222164 339276 222216
rect 299480 222096 299532 222148
rect 300768 222096 300820 222148
rect 298928 221552 298980 221604
rect 313372 221552 313424 221604
rect 57244 221484 57296 221536
rect 253388 221484 253440 221536
rect 297364 221484 297416 221536
rect 337384 221484 337436 221536
rect 59820 221416 59872 221468
rect 352288 221416 352340 221468
rect 226064 220804 226116 220856
rect 300768 220804 300820 220856
rect 578884 220804 578936 220856
rect 299020 220260 299072 220312
rect 306380 220260 306432 220312
rect 57152 220192 57204 220244
rect 291936 220192 291988 220244
rect 298836 220192 298888 220244
rect 328460 220192 328512 220244
rect 60556 220124 60608 220176
rect 294604 220124 294656 220176
rect 297272 220124 297324 220176
rect 336924 220124 336976 220176
rect 3608 220056 3660 220108
rect 510804 220056 510856 220108
rect 351276 219376 351328 219428
rect 579896 219376 579948 219428
rect 57888 218764 57940 218816
rect 253204 218764 253256 218816
rect 57612 218696 57664 218748
rect 293224 218696 293276 218748
rect 222936 216656 222988 216708
rect 296812 216656 296864 216708
rect 247684 215296 247736 215348
rect 297732 215296 297784 215348
rect 57244 214548 57296 214600
rect 57520 214548 57572 214600
rect 246304 213936 246356 213988
rect 297732 213936 297784 213988
rect 222292 212984 222344 213036
rect 226064 212984 226116 213036
rect 243544 212508 243596 212560
rect 297732 212508 297784 212560
rect 242164 211148 242216 211200
rect 297732 211148 297784 211200
rect 239404 209788 239456 209840
rect 297732 209788 297784 209840
rect 238024 208360 238076 208412
rect 297732 208360 297784 208412
rect 232504 207000 232556 207052
rect 297732 207000 297784 207052
rect 418804 206932 418856 206984
rect 580172 206932 580224 206984
rect 229744 205640 229796 205692
rect 297732 205640 297784 205692
rect 223212 205572 223264 205624
rect 229836 205572 229888 205624
rect 287704 201492 287756 201544
rect 296812 201492 296864 201544
rect 51724 201424 51776 201476
rect 57336 201424 57388 201476
rect 228364 200132 228416 200184
rect 297732 200132 297784 200184
rect 225604 198704 225656 198756
rect 297732 198704 297784 198756
rect 224316 197344 224368 197396
rect 297732 197344 297784 197396
rect 50988 197276 51040 197328
rect 57336 197276 57388 197328
rect 224224 195984 224276 196036
rect 297732 195984 297784 196036
rect 223488 194556 223540 194608
rect 233976 194556 234028 194608
rect 250444 194556 250496 194608
rect 297732 194556 297784 194608
rect 235264 193196 235316 193248
rect 297732 193196 297784 193248
rect 229836 193128 229888 193180
rect 297548 193128 297600 193180
rect 552664 193128 552716 193180
rect 580172 193128 580224 193180
rect 50896 192448 50948 192500
rect 57244 192448 57296 192500
rect 223488 191836 223540 191888
rect 229928 191836 229980 191888
rect 233884 190476 233936 190528
rect 297732 190476 297784 190528
rect 222844 190408 222896 190460
rect 297548 190408 297600 190460
rect 222844 189048 222896 189100
rect 224960 189048 225012 189100
rect 50436 188980 50488 189032
rect 57336 188980 57388 189032
rect 223028 188980 223080 189032
rect 297732 188980 297784 189032
rect 222844 186328 222896 186380
rect 228456 186328 228508 186380
rect 222936 186260 222988 186312
rect 297732 186260 297784 186312
rect 51080 184832 51132 184884
rect 56692 184832 56744 184884
rect 233976 184832 234028 184884
rect 297732 184832 297784 184884
rect 222292 183744 222344 183796
rect 225788 183744 225840 183796
rect 229928 183472 229980 183524
rect 297732 183472 297784 183524
rect 224960 182112 225012 182164
rect 297732 182112 297784 182164
rect 51172 180752 51224 180804
rect 56692 180752 56744 180804
rect 228456 180752 228508 180804
rect 297732 180752 297784 180804
rect 225788 179324 225840 179376
rect 297732 179324 297784 179376
rect 223488 177964 223540 178016
rect 297732 177964 297784 178016
rect 477868 177352 477920 177404
rect 516140 177352 516192 177404
rect 358452 177284 358504 177336
rect 426440 177284 426492 177336
rect 478512 177284 478564 177336
rect 520280 177284 520332 177336
rect 50344 176604 50396 176656
rect 57336 176604 57388 176656
rect 222660 176604 222712 176656
rect 297732 176604 297784 176656
rect 222660 175176 222712 175228
rect 297732 175176 297784 175228
rect 48872 173340 48924 173392
rect 57244 173340 57296 173392
rect 222384 173136 222436 173188
rect 297732 173136 297784 173188
rect 222476 171096 222528 171148
rect 297732 171096 297784 171148
rect 222936 169736 222988 169788
rect 297732 169736 297784 169788
rect 49516 169668 49568 169720
rect 57336 169668 57388 169720
rect 223488 167016 223540 167068
rect 297732 167016 297784 167068
rect 409144 166948 409196 167000
rect 580172 166948 580224 167000
rect 223028 165588 223080 165640
rect 296812 165588 296864 165640
rect 222936 164228 222988 164280
rect 297732 164228 297784 164280
rect 223488 162868 223540 162920
rect 297732 162868 297784 162920
rect 229100 161440 229152 161492
rect 297732 161440 297784 161492
rect 54576 161372 54628 161424
rect 57060 161372 57112 161424
rect 231124 160080 231176 160132
rect 297732 160080 297784 160132
rect 228456 158720 228508 158772
rect 297732 158720 297784 158772
rect 225696 157360 225748 157412
rect 296812 157360 296864 157412
rect 53104 157292 53156 157344
rect 57060 157292 57112 157344
rect 222568 157088 222620 157140
rect 229100 157088 229152 157140
rect 229836 155932 229888 155984
rect 297732 155932 297784 155984
rect 222936 154572 222988 154624
rect 297732 154572 297784 154624
rect 222844 153212 222896 153264
rect 297732 153212 297784 153264
rect 54484 153144 54536 153196
rect 57336 153144 57388 153196
rect 536104 153144 536156 153196
rect 579804 153144 579856 153196
rect 236644 151784 236696 151836
rect 297732 151784 297784 151836
rect 223488 150424 223540 150476
rect 231124 150424 231176 150476
rect 235356 149064 235408 149116
rect 297732 149064 297784 149116
rect 50804 148996 50856 149048
rect 57336 148996 57388 149048
rect 233976 147636 234028 147688
rect 296812 147636 296864 147688
rect 223488 147228 223540 147280
rect 228456 147228 228508 147280
rect 231124 146276 231176 146328
rect 297732 146276 297784 146328
rect 228456 144916 228508 144968
rect 297732 144916 297784 144968
rect 50712 144508 50764 144560
rect 57336 144508 57388 144560
rect 222476 144304 222528 144356
rect 225696 144304 225748 144356
rect 232596 143556 232648 143608
rect 297732 143556 297784 143608
rect 251824 142128 251876 142180
rect 297548 142128 297600 142180
rect 257344 142060 257396 142112
rect 297732 142060 297784 142112
rect 223488 141448 223540 141500
rect 229836 141448 229888 141500
rect 51264 140700 51316 140752
rect 57428 140700 57480 140752
rect 273996 140700 274048 140752
rect 297732 140700 297784 140752
rect 271236 139340 271288 139392
rect 297732 139340 297784 139392
rect 353944 139340 353996 139392
rect 580172 139340 580224 139392
rect 278044 137912 278096 137964
rect 297732 137912 297784 137964
rect 3148 137708 3200 137760
rect 8944 137708 8996 137760
rect 222476 137232 222528 137284
rect 236644 137232 236696 137284
rect 269856 136552 269908 136604
rect 296812 136552 296864 136604
rect 275376 135192 275428 135244
rect 297732 135192 297784 135244
rect 223120 133152 223172 133204
rect 235356 133152 235408 133204
rect 274088 132404 274140 132456
rect 297732 132404 297784 132456
rect 271328 131044 271380 131096
rect 297732 131044 297784 131096
rect 223488 130364 223540 130416
rect 233976 130364 234028 130416
rect 275468 129684 275520 129736
rect 297732 129684 297784 129736
rect 222476 128256 222528 128308
rect 231124 128256 231176 128308
rect 257436 128256 257488 128308
rect 297732 128256 297784 128308
rect 261576 126896 261628 126948
rect 297732 126896 297784 126948
rect 372896 126896 372948 126948
rect 580172 126896 580224 126948
rect 279424 125536 279476 125588
rect 297732 125536 297784 125588
rect 223212 124584 223264 124636
rect 228456 124584 228508 124636
rect 268476 124108 268528 124160
rect 297732 124108 297784 124160
rect 265716 122748 265768 122800
rect 297732 122748 297784 122800
rect 264336 121388 264388 121440
rect 297732 121388 297784 121440
rect 289084 120028 289136 120080
rect 297732 120028 297784 120080
rect 223488 118600 223540 118652
rect 232596 118600 232648 118652
rect 269948 118600 270000 118652
rect 296812 118600 296864 118652
rect 284944 117240 284996 117292
rect 297732 117240 297784 117292
rect 342904 117240 342956 117292
rect 475568 117240 475620 117292
rect 223488 115880 223540 115932
rect 251824 115880 251876 115932
rect 278228 114452 278280 114504
rect 297732 114452 297784 114504
rect 257528 113092 257580 113144
rect 297732 113092 297784 113144
rect 571984 113092 572036 113144
rect 580172 113092 580224 113144
rect 222200 112956 222252 113008
rect 224408 112956 224460 113008
rect 223488 110372 223540 110424
rect 247684 110372 247736 110424
rect 342904 108944 342956 108996
rect 481088 108944 481140 108996
rect 222660 107584 222712 107636
rect 246304 107584 246356 107636
rect 342904 106224 342956 106276
rect 505100 106224 505152 106276
rect 222844 104796 222896 104848
rect 243544 104796 243596 104848
rect 223488 102076 223540 102128
rect 242164 102076 242216 102128
rect 223028 99288 223080 99340
rect 239404 99288 239456 99340
rect 223120 96568 223172 96620
rect 238024 96568 238076 96620
rect 223488 93780 223540 93832
rect 232504 93780 232556 93832
rect 223396 91740 223448 91792
rect 295984 91740 296036 91792
rect 223488 90312 223540 90364
rect 229744 90312 229796 90364
rect 264244 90312 264296 90364
rect 296812 90312 296864 90364
rect 358544 89020 358596 89072
rect 408500 89020 408552 89072
rect 260196 88952 260248 89004
rect 297364 88952 297416 89004
rect 358636 88952 358688 89004
rect 415400 88952 415452 89004
rect 340420 88680 340472 88732
rect 342536 88680 342588 88732
rect 291844 88272 291896 88324
rect 298008 88272 298060 88324
rect 223488 87592 223540 87644
rect 287704 87592 287756 87644
rect 358820 86912 358872 86964
rect 580172 86912 580224 86964
rect 3148 85484 3200 85536
rect 14464 85484 14516 85536
rect 267004 85484 267056 85536
rect 297548 85484 297600 85536
rect 269764 84124 269816 84176
rect 297916 84124 297968 84176
rect 275284 82764 275336 82816
rect 297916 82764 297968 82816
rect 223488 81336 223540 81388
rect 228364 81336 228416 81388
rect 273904 79976 273956 80028
rect 298008 79976 298060 80028
rect 271144 78616 271196 78668
rect 297548 78616 297600 78668
rect 222476 78548 222528 78600
rect 225604 78548 225656 78600
rect 260104 77188 260156 77240
rect 297180 77188 297232 77240
rect 255964 75828 256016 75880
rect 298008 75828 298060 75880
rect 222200 75692 222252 75744
rect 224316 75692 224368 75744
rect 261484 74468 261536 74520
rect 298008 74468 298060 74520
rect 256056 73108 256108 73160
rect 296812 73108 296864 73160
rect 480996 73108 481048 73160
rect 580172 73108 580224 73160
rect 222200 73040 222252 73092
rect 224224 73040 224276 73092
rect 223488 70320 223540 70372
rect 250444 70320 250496 70372
rect 265624 70320 265676 70372
rect 298008 70320 298060 70372
rect 343088 69028 343140 69080
rect 489920 69028 489972 69080
rect 268384 68960 268436 69012
rect 297180 68960 297232 69012
rect 223488 67532 223540 67584
rect 235264 67532 235316 67584
rect 282184 67532 282236 67584
rect 297548 67532 297600 67584
rect 343180 66240 343232 66292
rect 482376 66240 482428 66292
rect 222844 64812 222896 64864
rect 233884 64812 233936 64864
rect 278136 64812 278188 64864
rect 297916 64812 297968 64864
rect 343180 63520 343232 63572
rect 418804 63520 418856 63572
rect 342352 62704 342404 62756
rect 343180 62704 343232 62756
rect 342352 62092 342404 62144
rect 480352 62092 480404 62144
rect 264428 62024 264480 62076
rect 298008 62024 298060 62076
rect 215300 61548 215352 61600
rect 342720 61548 342772 61600
rect 168380 61480 168432 61532
rect 341708 61480 341760 61532
rect 158720 61412 158772 61464
rect 343088 61412 343140 61464
rect 154580 61344 154632 61396
rect 342996 61344 343048 61396
rect 356704 60664 356756 60716
rect 580172 60664 580224 60716
rect 296628 60188 296680 60240
rect 303620 60188 303672 60240
rect 295248 60120 295300 60172
rect 310520 60120 310572 60172
rect 314660 60120 314712 60172
rect 352564 60120 352616 60172
rect 211160 60052 211212 60104
rect 342812 60052 342864 60104
rect 193220 59984 193272 60036
rect 341340 59984 341392 60036
rect 3056 59304 3108 59356
rect 369124 59304 369176 59356
rect 172520 58692 172572 58744
rect 341616 58692 341668 58744
rect 133880 58624 133932 58676
rect 340512 58624 340564 58676
rect 229100 57332 229152 57384
rect 342444 57332 342496 57384
rect 190460 57264 190512 57316
rect 340328 57264 340380 57316
rect 176660 57196 176712 57248
rect 341524 57196 341576 57248
rect 233240 55972 233292 56024
rect 343180 55972 343232 56024
rect 226340 55904 226392 55956
rect 341248 55904 341300 55956
rect 179420 55836 179472 55888
rect 341432 55836 341484 55888
rect 247040 54612 247092 54664
rect 340144 54612 340196 54664
rect 218060 54544 218112 54596
rect 342628 54544 342680 54596
rect 204260 54476 204312 54528
rect 340236 54476 340288 54528
rect 346400 53048 346452 53100
rect 509792 53048 509844 53100
rect 251180 50328 251232 50380
rect 341064 50328 341116 50380
rect 201500 47540 201552 47592
rect 491944 47540 491996 47592
rect 359556 46860 359608 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 472716 45500 472768 45552
rect 99380 43392 99432 43444
rect 513012 43392 513064 43444
rect 151820 42032 151872 42084
rect 342904 42032 342956 42084
rect 208400 40808 208452 40860
rect 341156 40808 341208 40860
rect 120080 40740 120132 40792
rect 481272 40740 481324 40792
rect 56600 40672 56652 40724
rect 512276 40672 512328 40724
rect 113180 37884 113232 37936
rect 462964 37884 463016 37936
rect 117320 36524 117372 36576
rect 436744 36524 436796 36576
rect 236000 35300 236052 35352
rect 340052 35300 340104 35352
rect 110420 35232 110472 35284
rect 496176 35232 496228 35284
rect 23480 35164 23532 35216
rect 416044 35164 416096 35216
rect 70400 33736 70452 33788
rect 501236 33736 501288 33788
rect 480904 33056 480956 33108
rect 580172 33056 580224 33108
rect 378140 31016 378192 31068
rect 476856 31016 476908 31068
rect 77300 29588 77352 29640
rect 502984 29588 503036 29640
rect 92480 26868 92532 26920
rect 493416 26868 493468 26920
rect 371240 22720 371292 22772
rect 440884 22720 440936 22772
rect 396172 21428 396224 21480
rect 422944 21428 422996 21480
rect 423772 21428 423824 21480
rect 504456 21428 504508 21480
rect 60740 21360 60792 21412
rect 475476 21360 475528 21412
rect 3424 20612 3476 20664
rect 510712 20612 510764 20664
rect 102140 19932 102192 19984
rect 496084 19932 496136 19984
rect 197360 18708 197412 18760
rect 340972 18708 341024 18760
rect 360200 18708 360252 18760
rect 450544 18708 450596 18760
rect 106280 18640 106332 18692
rect 405004 18640 405056 18692
rect 19340 18572 19392 18624
rect 402244 18572 402296 18624
rect 420184 17280 420236 17332
rect 498292 17280 498344 17332
rect 357440 17212 357492 17264
rect 454684 17212 454736 17264
rect 390928 15920 390980 15972
rect 440240 15920 440292 15972
rect 81624 15852 81676 15904
rect 493324 15852 493376 15904
rect 254216 14424 254268 14476
rect 494796 14424 494848 14476
rect 353576 13064 353628 13116
rect 476764 13064 476816 13116
rect 378692 11704 378744 11756
rect 455696 11704 455748 11756
rect 242900 10344 242952 10396
rect 342260 10344 342312 10396
rect 240140 10276 240192 10328
rect 340880 10276 340932 10328
rect 477868 10276 477920 10328
rect 494704 10276 494756 10328
rect 445024 9052 445076 9104
rect 494704 9052 494756 9104
rect 89168 8984 89220 9036
rect 510344 8984 510396 9036
rect 85672 8916 85724 8968
rect 509976 8916 510028 8968
rect 396080 8236 396132 8288
rect 402520 8236 402572 8288
rect 482376 8236 482428 8288
rect 487620 8236 487672 8288
rect 418804 7760 418856 7812
rect 484032 7760 484084 7812
rect 67916 7692 67968 7744
rect 475384 7692 475436 7744
rect 478696 7692 478748 7744
rect 581000 7692 581052 7744
rect 64328 7624 64380 7676
rect 512828 7624 512880 7676
rect 4068 7556 4120 7608
rect 510620 7556 510672 7608
rect 359464 6808 359516 6860
rect 580172 6808 580224 6860
rect 46664 6264 46716 6316
rect 489644 6264 489696 6316
rect 35992 6196 36044 6248
rect 491576 6196 491628 6248
rect 39580 6128 39632 6180
rect 499948 6128 500000 6180
rect 141240 4972 141292 5024
rect 357624 4972 357676 5024
rect 473452 4972 473504 5024
rect 477960 4972 478012 5024
rect 559748 4972 559800 5024
rect 342536 4904 342588 4956
rect 350448 4904 350500 4956
rect 508320 4904 508372 4956
rect 50160 4836 50212 4888
rect 507676 4836 507728 4888
rect 2872 4768 2924 4820
rect 512736 4768 512788 4820
rect 339868 3952 339920 4004
rect 353392 3952 353444 4004
rect 332692 3884 332744 3936
rect 350540 3884 350592 3936
rect 336280 3816 336332 3868
rect 355416 3816 355468 3868
rect 296536 3748 296588 3800
rect 322112 3748 322164 3800
rect 325608 3748 325660 3800
rect 351184 3748 351236 3800
rect 307944 3680 307996 3732
rect 355324 3680 355376 3732
rect 538864 3680 538916 3732
rect 556160 3680 556212 3732
rect 222752 3612 222804 3664
rect 340420 3612 340472 3664
rect 343364 3612 343416 3664
rect 353300 3612 353352 3664
rect 453304 3612 453356 3664
rect 508504 3612 508556 3664
rect 530584 3612 530636 3664
rect 102140 3544 102192 3596
rect 103336 3544 103388 3596
rect 124680 3544 124732 3596
rect 489000 3544 489052 3596
rect 526444 3544 526496 3596
rect 531320 3544 531372 3596
rect 531964 3612 532016 3664
rect 541992 3612 542044 3664
rect 538404 3544 538456 3596
rect 544384 3544 544436 3596
rect 573916 3544 573968 3596
rect 32404 3476 32456 3528
rect 472624 3476 472676 3528
rect 479432 3476 479484 3528
rect 485228 3476 485280 3528
rect 498200 3476 498252 3528
rect 499028 3476 499080 3528
rect 522304 3476 522356 3528
rect 524236 3476 524288 3528
rect 525064 3476 525116 3528
rect 527824 3476 527876 3528
rect 534724 3476 534776 3528
rect 28908 3408 28960 3460
rect 468484 3408 468536 3460
rect 482284 3408 482336 3460
rect 510068 3408 510120 3460
rect 527916 3408 527968 3460
rect 534908 3408 534960 3460
rect 549904 3476 549956 3528
rect 545488 3408 545540 3460
rect 545764 3408 545816 3460
rect 577412 3408 577464 3460
rect 578884 3476 578936 3528
rect 579804 3476 579856 3528
rect 582196 3408 582248 3460
rect 143540 3340 143592 3392
rect 144736 3340 144788 3392
rect 168380 3340 168432 3392
rect 169576 3340 169628 3392
rect 193220 3340 193272 3392
rect 194416 3340 194468 3392
rect 218060 3340 218112 3392
rect 219256 3340 219308 3392
rect 242900 3340 242952 3392
rect 244096 3340 244148 3392
rect 414664 3340 414716 3392
rect 420184 3340 420236 3392
rect 423772 3340 423824 3392
rect 424968 3340 425020 3392
rect 448520 3340 448572 3392
rect 449808 3340 449860 3392
rect 398840 3136 398892 3188
rect 400128 3136 400180 3188
rect 415400 3136 415452 3188
rect 416688 3136 416740 3188
rect 440240 3136 440292 3188
rect 441528 3136 441580 3188
rect 506480 3136 506532 3188
rect 508964 3136 509016 3188
rect 374000 3000 374052 3052
rect 375288 3000 375340 3052
<< metal2 >>
rect 6932 703582 7972 703610
rect 6932 665854 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700330 24348 703520
rect 72988 700398 73016 703520
rect 89180 700466 89208 703520
rect 89168 700460 89220 700466
rect 89168 700402 89220 700408
rect 72976 700392 73028 700398
rect 72976 700334 73028 700340
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 105464 697610 105492 703520
rect 105452 697604 105504 697610
rect 105452 697546 105504 697552
rect 6920 665848 6972 665854
rect 6920 665790 6972 665796
rect 52092 663876 52144 663882
rect 52092 663818 52144 663824
rect 46480 663808 46532 663814
rect 46480 663750 46532 663756
rect 3698 662688 3754 662697
rect 3698 662623 3754 662632
rect 45468 662652 45520 662658
rect 3514 662552 3570 662561
rect 3514 662487 3570 662496
rect 3424 661156 3476 661162
rect 3424 661098 3476 661104
rect 3332 659864 3384 659870
rect 3332 659806 3384 659812
rect 3344 658209 3372 659806
rect 3330 658200 3386 658209
rect 3330 658135 3386 658144
rect 3436 449585 3464 661098
rect 3528 462641 3556 662487
rect 3608 661224 3660 661230
rect 3608 661166 3660 661172
rect 3620 501809 3648 661166
rect 3712 514865 3740 662623
rect 45468 662594 45520 662600
rect 3792 661088 3844 661094
rect 3792 661030 3844 661036
rect 3804 553897 3832 661030
rect 3790 553888 3846 553897
rect 3790 553823 3846 553832
rect 3698 514856 3754 514865
rect 3698 514791 3754 514800
rect 3606 501800 3662 501809
rect 3606 501735 3662 501744
rect 45480 467838 45508 662594
rect 46388 662448 46440 662454
rect 46388 662390 46440 662396
rect 46400 473346 46428 662390
rect 46388 473340 46440 473346
rect 46388 473282 46440 473288
rect 45468 467832 45520 467838
rect 45468 467774 45520 467780
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 46492 456414 46520 663750
rect 50986 663232 51042 663241
rect 50986 663167 51042 663176
rect 50436 663128 50488 663134
rect 46570 663096 46626 663105
rect 50436 663070 50488 663076
rect 46570 663031 46626 663040
rect 46756 663060 46808 663066
rect 46480 456408 46532 456414
rect 46480 456350 46532 456356
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 46584 445738 46612 663031
rect 46756 663002 46808 663008
rect 46662 662960 46718 662969
rect 46662 662895 46718 662904
rect 46572 445732 46624 445738
rect 46572 445674 46624 445680
rect 46676 438870 46704 662895
rect 46664 438864 46716 438870
rect 46664 438806 46716 438812
rect 46768 433294 46796 663002
rect 47860 662720 47912 662726
rect 47860 662662 47912 662668
rect 46848 660068 46900 660074
rect 46848 660010 46900 660016
rect 46756 433288 46808 433294
rect 46756 433230 46808 433236
rect 46860 427786 46888 660010
rect 47872 462330 47900 662662
rect 50066 661872 50122 661881
rect 50066 661807 50122 661816
rect 49974 661736 50030 661745
rect 49974 661671 50030 661680
rect 49330 661600 49386 661609
rect 49148 661564 49200 661570
rect 49330 661535 49386 661544
rect 49148 661506 49200 661512
rect 48962 661464 49018 661473
rect 48962 661399 49018 661408
rect 48870 661056 48926 661065
rect 48870 660991 48926 661000
rect 48134 660648 48190 660657
rect 48134 660583 48190 660592
rect 48042 660512 48098 660521
rect 48042 660447 48098 660456
rect 47950 660376 48006 660385
rect 47950 660311 48006 660320
rect 47860 462324 47912 462330
rect 47860 462266 47912 462272
rect 46848 427780 46900 427786
rect 46848 427722 46900 427728
rect 47964 421297 47992 660311
rect 47950 421288 48006 421297
rect 47950 421223 48006 421232
rect 48056 415449 48084 660447
rect 48042 415440 48098 415449
rect 48042 415375 48098 415384
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 48148 409601 48176 660583
rect 48594 660240 48650 660249
rect 48594 660175 48650 660184
rect 48228 660136 48280 660142
rect 48228 660078 48280 660084
rect 48134 409592 48190 409601
rect 48134 409527 48190 409536
rect 48240 403753 48268 660078
rect 48608 585041 48636 660175
rect 48778 659968 48834 659977
rect 48778 659903 48834 659912
rect 48688 652792 48740 652798
rect 48688 652734 48740 652740
rect 48594 585032 48650 585041
rect 48594 584967 48650 584976
rect 48700 579193 48728 652734
rect 48792 620129 48820 659903
rect 48778 620120 48834 620129
rect 48778 620055 48834 620064
rect 48780 619064 48832 619070
rect 48780 619006 48832 619012
rect 48686 579184 48742 579193
rect 48686 579119 48742 579128
rect 48792 555801 48820 619006
rect 48884 596737 48912 660991
rect 48870 596728 48926 596737
rect 48870 596663 48926 596672
rect 48976 590889 49004 661399
rect 49056 641776 49108 641782
rect 49056 641718 49108 641724
rect 48962 590880 49018 590889
rect 48962 590815 49018 590824
rect 49068 567497 49096 641718
rect 49160 631825 49188 661506
rect 49240 660204 49292 660210
rect 49240 660146 49292 660152
rect 49252 649369 49280 660146
rect 49238 649360 49294 649369
rect 49238 649295 49294 649304
rect 49240 648576 49292 648582
rect 49240 648518 49292 648524
rect 49146 631816 49202 631825
rect 49146 631751 49202 631760
rect 49148 629400 49200 629406
rect 49148 629342 49200 629348
rect 49054 567488 49110 567497
rect 49054 567423 49110 567432
rect 48778 555792 48834 555801
rect 48778 555727 48834 555736
rect 49160 549953 49188 629342
rect 49252 561649 49280 648518
rect 49344 573345 49372 661535
rect 49792 661292 49844 661298
rect 49792 661234 49844 661240
rect 49424 660612 49476 660618
rect 49424 660554 49476 660560
rect 49436 637673 49464 660554
rect 49608 660544 49660 660550
rect 49608 660486 49660 660492
rect 49516 660272 49568 660278
rect 49516 660214 49568 660220
rect 49528 654134 49556 660214
rect 49620 655217 49648 660486
rect 49804 659705 49832 661234
rect 49790 659696 49846 659705
rect 49790 659631 49846 659640
rect 49606 655208 49662 655217
rect 49606 655143 49662 655152
rect 49528 654106 49648 654134
rect 49620 643521 49648 654106
rect 49988 652798 50016 661671
rect 50080 658050 50108 661807
rect 50252 661768 50304 661774
rect 50252 661710 50304 661716
rect 50160 660476 50212 660482
rect 50160 660418 50212 660424
rect 50172 659841 50200 660418
rect 50158 659832 50214 659841
rect 50158 659767 50214 659776
rect 50080 658022 50200 658050
rect 49976 652792 50028 652798
rect 49976 652734 50028 652740
rect 50172 648582 50200 658022
rect 50160 648576 50212 648582
rect 50160 648518 50212 648524
rect 49606 643512 49662 643521
rect 49606 643447 49662 643456
rect 50264 641782 50292 661710
rect 50344 660340 50396 660346
rect 50344 660282 50396 660288
rect 50356 659705 50384 660282
rect 50342 659696 50398 659705
rect 50342 659631 50398 659640
rect 50344 658708 50396 658714
rect 50344 658650 50396 658656
rect 50252 641776 50304 641782
rect 50252 641718 50304 641724
rect 49422 637664 49478 637673
rect 49422 637599 49478 637608
rect 49424 636744 49476 636750
rect 49424 636686 49476 636692
rect 49330 573336 49386 573345
rect 49330 573271 49386 573280
rect 49238 561640 49294 561649
rect 49238 561575 49294 561584
rect 49146 549944 49202 549953
rect 49146 549879 49202 549888
rect 49436 544105 49464 636686
rect 50356 619070 50384 658650
rect 50448 629406 50476 663070
rect 50896 662856 50948 662862
rect 50896 662798 50948 662804
rect 50528 661632 50580 661638
rect 50528 661574 50580 661580
rect 50540 636750 50568 661574
rect 50804 661496 50856 661502
rect 50804 661438 50856 661444
rect 50620 661428 50672 661434
rect 50620 661370 50672 661376
rect 50528 636744 50580 636750
rect 50528 636686 50580 636692
rect 50436 629400 50488 629406
rect 50436 629342 50488 629348
rect 50344 619064 50396 619070
rect 50344 619006 50396 619012
rect 49516 594856 49568 594862
rect 49516 594798 49568 594804
rect 49422 544096 49478 544105
rect 49422 544031 49478 544040
rect 49422 539608 49478 539617
rect 49422 539543 49478 539552
rect 49436 538257 49464 539543
rect 49422 538248 49478 538257
rect 49422 538183 49478 538192
rect 49330 521656 49386 521665
rect 49330 521591 49386 521600
rect 49344 520713 49372 521591
rect 49330 520704 49386 520713
rect 49330 520639 49386 520648
rect 49238 503160 49294 503169
rect 49238 503095 49294 503104
rect 48870 496904 48926 496913
rect 48870 496839 48926 496848
rect 48778 468072 48834 468081
rect 48778 468007 48834 468016
rect 48792 467838 48820 468007
rect 48780 467832 48832 467838
rect 48780 467774 48832 467780
rect 48320 445732 48372 445738
rect 48320 445674 48372 445680
rect 48332 444689 48360 445674
rect 48318 444680 48374 444689
rect 48318 444615 48374 444624
rect 48320 438864 48372 438870
rect 48318 438832 48320 438841
rect 48372 438832 48374 438841
rect 48318 438767 48374 438776
rect 48226 403744 48282 403753
rect 48226 403679 48282 403688
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3436 281518 3464 397423
rect 48318 392048 48374 392057
rect 46848 392012 46900 392018
rect 48318 391983 48320 391992
rect 46848 391954 46900 391960
rect 48372 391983 48374 391992
rect 48320 391954 48372 391960
rect 46756 385076 46808 385082
rect 46756 385018 46808 385024
rect 46664 379568 46716 379574
rect 46664 379510 46716 379516
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 282062 3556 306167
rect 3606 293176 3662 293185
rect 3606 293111 3662 293120
rect 3516 282056 3568 282062
rect 3516 281998 3568 282004
rect 3424 281512 3476 281518
rect 3424 281454 3476 281460
rect 3620 280090 3648 293111
rect 3608 280084 3660 280090
rect 3608 280026 3660 280032
rect 46676 280022 46704 379510
rect 46768 281926 46796 385018
rect 46756 281920 46808 281926
rect 46756 281862 46808 281868
rect 46664 280016 46716 280022
rect 46664 279958 46716 279964
rect 46860 279954 46888 391954
rect 48318 386200 48374 386209
rect 48318 386135 48374 386144
rect 48332 385082 48360 386135
rect 48320 385076 48372 385082
rect 48320 385018 48372 385024
rect 48226 374504 48282 374513
rect 48226 374439 48282 374448
rect 48134 368656 48190 368665
rect 48134 368591 48190 368600
rect 48042 362808 48098 362817
rect 48042 362743 48098 362752
rect 47950 351112 48006 351121
rect 47950 351047 48006 351056
rect 47858 345264 47914 345273
rect 47858 345199 47914 345208
rect 47872 281217 47900 345199
rect 47964 281353 47992 351047
rect 47950 281344 48006 281353
rect 47950 281279 48006 281288
rect 47858 281208 47914 281217
rect 47858 281143 47914 281152
rect 48056 280974 48084 362743
rect 48044 280968 48096 280974
rect 48044 280910 48096 280916
rect 48148 280537 48176 368591
rect 48134 280528 48190 280537
rect 48134 280463 48190 280472
rect 46848 279948 46900 279954
rect 46848 279890 46900 279896
rect 48240 279886 48268 374439
rect 48686 298480 48742 298489
rect 48686 298415 48742 298424
rect 48700 281110 48728 298415
rect 48778 292632 48834 292641
rect 48778 292567 48834 292576
rect 48792 281858 48820 292567
rect 48780 281852 48832 281858
rect 48780 281794 48832 281800
rect 48688 281104 48740 281110
rect 48688 281046 48740 281052
rect 48228 279880 48280 279886
rect 48228 279822 48280 279828
rect 8944 276684 8996 276690
rect 8944 276626 8996 276632
rect 3424 268388 3476 268394
rect 3424 268330 3476 268336
rect 3436 254153 3464 268330
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3424 241460 3476 241466
rect 3424 241402 3476 241408
rect 3436 241097 3464 241402
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3516 225616 3568 225622
rect 3516 225558 3568 225564
rect 3424 224324 3476 224330
rect 3424 224266 3476 224272
rect 3148 137760 3200 137766
rect 3148 137702 3200 137708
rect 3160 136785 3188 137702
rect 3146 136776 3202 136785
rect 3146 136711 3202 136720
rect 3436 97617 3464 224266
rect 3528 149841 3556 225558
rect 3700 224256 3752 224262
rect 3700 224198 3752 224204
rect 3608 220108 3660 220114
rect 3608 220050 3660 220056
rect 3620 188873 3648 220050
rect 3712 201929 3740 224198
rect 3698 201920 3754 201929
rect 3698 201855 3754 201864
rect 3606 188864 3662 188873
rect 3606 188799 3662 188808
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 8956 137766 8984 276626
rect 13820 268456 13872 268462
rect 13820 268398 13872 268404
rect 9680 239420 9732 239426
rect 9680 239362 9732 239368
rect 8944 137760 8996 137766
rect 8944 137702 8996 137708
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 4080 6497 4108 7550
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2884 480 2912 4762
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 239362
rect 13832 16574 13860 268398
rect 14464 233912 14516 233918
rect 14464 233854 14516 233860
rect 14476 85542 14504 233854
rect 42800 225684 42852 225690
rect 42800 225626 42852 225632
rect 14464 85536 14516 85542
rect 14464 85478 14516 85484
rect 23480 35216 23532 35222
rect 23480 35158 23532 35164
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19352 16574 19380 18566
rect 23492 16574 23520 35158
rect 13832 16546 14320 16574
rect 19352 16546 19472 16574
rect 23492 16546 24256 16574
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 19444 480 19472 16546
rect 24228 480 24256 16546
rect 35992 6248 36044 6254
rect 35992 6190 36044 6196
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 28908 3460 28960 3466
rect 28908 3402 28960 3408
rect 28920 480 28948 3402
rect 32416 480 32444 3470
rect 36004 480 36032 6190
rect 39580 6180 39632 6186
rect 39580 6122 39632 6128
rect 39592 480 39620 6122
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42812 354 42840 225626
rect 48884 173398 48912 496839
rect 49252 495514 49280 503095
rect 49240 495508 49292 495514
rect 49240 495450 49292 495456
rect 49344 481642 49372 520639
rect 49436 485858 49464 538183
rect 49528 491473 49556 594798
rect 49608 590640 49660 590646
rect 49608 590582 49660 590588
rect 49620 497321 49648 590582
rect 49606 497312 49662 497321
rect 49606 497247 49662 497256
rect 49620 496913 49648 497247
rect 49606 496904 49662 496913
rect 49606 496839 49662 496848
rect 50344 495508 50396 495514
rect 50344 495450 50396 495456
rect 49514 491464 49570 491473
rect 49514 491399 49570 491408
rect 49424 485852 49476 485858
rect 49424 485794 49476 485800
rect 49332 481636 49384 481642
rect 49332 481578 49384 481584
rect 48962 473920 49018 473929
rect 48962 473855 49018 473864
rect 48976 473346 49004 473855
rect 48964 473340 49016 473346
rect 48964 473282 49016 473288
rect 48976 281314 49004 473282
rect 49056 467832 49108 467838
rect 49056 467774 49108 467780
rect 48964 281308 49016 281314
rect 48964 281250 49016 281256
rect 49068 281178 49096 467774
rect 49148 433288 49200 433294
rect 49148 433230 49200 433236
rect 49160 432993 49188 433230
rect 49146 432984 49202 432993
rect 49146 432919 49202 432928
rect 49424 427780 49476 427786
rect 49424 427722 49476 427728
rect 49436 427145 49464 427722
rect 49422 427136 49478 427145
rect 49422 427071 49478 427080
rect 49422 380352 49478 380361
rect 49422 380287 49478 380296
rect 49436 379574 49464 380287
rect 49424 379568 49476 379574
rect 49424 379510 49476 379516
rect 49422 327720 49478 327729
rect 49422 327655 49478 327664
rect 49330 321872 49386 321881
rect 49330 321807 49386 321816
rect 49238 316024 49294 316033
rect 49238 315959 49294 315968
rect 49146 304328 49202 304337
rect 49146 304263 49202 304272
rect 49160 281382 49188 304263
rect 49148 281376 49200 281382
rect 49148 281318 49200 281324
rect 49056 281172 49108 281178
rect 49056 281114 49108 281120
rect 49252 281042 49280 315959
rect 49240 281036 49292 281042
rect 49240 280978 49292 280984
rect 49344 280945 49372 321807
rect 49436 281081 49464 327655
rect 49422 281072 49478 281081
rect 49422 281007 49478 281016
rect 49330 280936 49386 280945
rect 49330 280871 49386 280880
rect 48872 173392 48924 173398
rect 48872 173334 48924 173340
rect 49528 169726 49556 491399
rect 49792 456408 49844 456414
rect 49790 456376 49792 456385
rect 49844 456376 49846 456385
rect 49790 456311 49846 456320
rect 50252 345092 50304 345098
rect 50252 345034 50304 345040
rect 50264 280158 50292 345034
rect 50252 280152 50304 280158
rect 50252 280094 50304 280100
rect 50356 176662 50384 495450
rect 50436 481636 50488 481642
rect 50436 481578 50488 481584
rect 50448 189038 50476 481578
rect 50632 450770 50660 661370
rect 50712 660408 50764 660414
rect 50712 660350 50764 660356
rect 50724 625977 50752 660350
rect 50710 625968 50766 625977
rect 50710 625903 50766 625912
rect 50816 509017 50844 661438
rect 50908 526561 50936 662798
rect 51000 658714 51028 663167
rect 51724 662992 51776 662998
rect 51724 662934 51776 662940
rect 51080 662924 51132 662930
rect 51080 662866 51132 662872
rect 50988 658708 51040 658714
rect 50988 658650 51040 658656
rect 50988 651432 51040 651438
rect 50988 651374 51040 651380
rect 51000 532409 51028 651374
rect 50986 532400 51042 532409
rect 50986 532335 51042 532344
rect 50894 526552 50950 526561
rect 50894 526487 50950 526496
rect 50802 509008 50858 509017
rect 50802 508943 50858 508952
rect 50816 507890 50844 508943
rect 50804 507884 50856 507890
rect 50804 507826 50856 507832
rect 50804 462324 50856 462330
rect 50804 462266 50856 462272
rect 50816 462233 50844 462266
rect 50802 462224 50858 462233
rect 50802 462159 50858 462168
rect 50710 456376 50766 456385
rect 50710 456311 50766 456320
rect 50620 450764 50672 450770
rect 50620 450706 50672 450712
rect 50528 409896 50580 409902
rect 50528 409838 50580 409844
rect 50540 281450 50568 409838
rect 50620 357468 50672 357474
rect 50620 357410 50672 357416
rect 50632 281994 50660 357410
rect 50620 281988 50672 281994
rect 50620 281930 50672 281936
rect 50528 281444 50580 281450
rect 50528 281386 50580 281392
rect 50436 189032 50488 189038
rect 50436 188974 50488 188980
rect 50344 176656 50396 176662
rect 50344 176598 50396 176604
rect 49516 169720 49568 169726
rect 49516 169662 49568 169668
rect 50724 144566 50752 456311
rect 50816 149054 50844 462159
rect 50908 192506 50936 526487
rect 51000 197334 51028 532335
rect 51092 514865 51120 662866
rect 51170 662824 51226 662833
rect 51170 662759 51226 662768
rect 51184 654134 51212 662759
rect 51356 660000 51408 660006
rect 51356 659942 51408 659948
rect 51264 659932 51316 659938
rect 51264 659874 51316 659880
rect 51276 659705 51304 659874
rect 51262 659696 51318 659705
rect 51262 659631 51318 659640
rect 51184 654106 51304 654134
rect 51078 514856 51134 514865
rect 51078 514791 51134 514800
rect 50988 197328 51040 197334
rect 50988 197270 51040 197276
rect 50896 192500 50948 192506
rect 50896 192442 50948 192448
rect 51092 184890 51120 514791
rect 51172 507884 51224 507890
rect 51172 507826 51224 507832
rect 51080 184884 51132 184890
rect 51080 184826 51132 184832
rect 51184 180810 51212 507826
rect 51276 485625 51304 654106
rect 51262 485616 51318 485625
rect 51262 485551 51318 485560
rect 51276 484401 51304 485551
rect 51262 484392 51318 484401
rect 51262 484327 51318 484336
rect 51264 450764 51316 450770
rect 51264 450706 51316 450712
rect 51276 450537 51304 450706
rect 51262 450528 51318 450537
rect 51262 450463 51318 450472
rect 51172 180804 51224 180810
rect 51172 180746 51224 180752
rect 50804 149048 50856 149054
rect 50804 148990 50856 148996
rect 50712 144560 50764 144566
rect 50712 144502 50764 144508
rect 51276 140758 51304 450463
rect 51368 397905 51396 659942
rect 51736 590646 51764 662934
rect 52000 662788 52052 662794
rect 52000 662730 52052 662736
rect 51908 662584 51960 662590
rect 51908 662526 51960 662532
rect 51816 661360 51868 661366
rect 51816 661302 51868 661308
rect 51828 594862 51856 661302
rect 51920 600817 51948 662526
rect 52012 607209 52040 662730
rect 52104 612785 52132 663818
rect 52184 662516 52236 662522
rect 52184 662458 52236 662464
rect 52196 651438 52224 662458
rect 136652 661706 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700534 154160 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 154120 700528 154172 700534
rect 154120 700470 154172 700476
rect 201512 661842 201540 702986
rect 218992 700602 219020 703520
rect 235184 700670 235212 703520
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 253296 700664 253348 700670
rect 253296 700606 253348 700612
rect 218980 700596 219032 700602
rect 218980 700538 219032 700544
rect 253204 700392 253256 700398
rect 253204 700334 253256 700340
rect 201500 661836 201552 661842
rect 201500 661778 201552 661784
rect 136640 661700 136692 661706
rect 136640 661642 136692 661648
rect 52184 651432 52236 651438
rect 52184 651374 52236 651380
rect 52090 612776 52146 612785
rect 52090 612711 52146 612720
rect 51998 607200 52054 607209
rect 51998 607135 52054 607144
rect 51906 600808 51962 600817
rect 51906 600743 51962 600752
rect 51816 594856 51868 594862
rect 51816 594798 51868 594804
rect 51724 590640 51776 590646
rect 51724 590582 51776 590588
rect 253216 555490 253244 700334
rect 253308 565146 253336 700606
rect 253388 700596 253440 700602
rect 253388 700538 253440 700544
rect 253400 569226 253428 700538
rect 264336 700528 264388 700534
rect 264336 700470 264388 700476
rect 257436 660612 257488 660618
rect 257436 660554 257488 660560
rect 254582 658200 254638 658209
rect 254582 658135 254638 658144
rect 254596 656946 254624 658135
rect 254584 656940 254636 656946
rect 254584 656882 254636 656888
rect 254582 652352 254638 652361
rect 254582 652287 254638 652296
rect 253938 646504 253994 646513
rect 253938 646439 253994 646448
rect 253952 645930 253980 646439
rect 253940 645924 253992 645930
rect 253940 645866 253992 645872
rect 254490 640656 254546 640665
rect 254490 640591 254546 640600
rect 254504 640354 254532 640591
rect 254492 640348 254544 640354
rect 254492 640290 254544 640296
rect 254398 634808 254454 634817
rect 254398 634743 254454 634752
rect 254412 633486 254440 634743
rect 254400 633480 254452 633486
rect 254400 633422 254452 633428
rect 254306 628960 254362 628969
rect 254306 628895 254362 628904
rect 254320 627978 254348 628895
rect 254308 627972 254360 627978
rect 254308 627914 254360 627920
rect 254030 623112 254086 623121
rect 254030 623047 254086 623056
rect 254044 622470 254072 623047
rect 254032 622464 254084 622470
rect 254032 622406 254084 622412
rect 254490 611416 254546 611425
rect 254490 611351 254492 611360
rect 254544 611351 254546 611360
rect 254492 611322 254544 611328
rect 254214 605568 254270 605577
rect 254214 605503 254270 605512
rect 254228 604518 254256 605503
rect 254216 604512 254268 604518
rect 254216 604454 254268 604460
rect 254122 599720 254178 599729
rect 254122 599655 254178 599664
rect 254136 599010 254164 599655
rect 254124 599004 254176 599010
rect 254124 598946 254176 598952
rect 254490 588024 254546 588033
rect 254490 587959 254492 587968
rect 254544 587959 254546 587968
rect 254492 587930 254544 587936
rect 253938 582176 253994 582185
rect 253938 582111 253994 582120
rect 253952 581330 253980 582111
rect 253940 581324 253992 581330
rect 253940 581266 253992 581272
rect 254490 576328 254546 576337
rect 254490 576263 254546 576272
rect 254504 575550 254532 576263
rect 254492 575544 254544 575550
rect 254492 575486 254544 575492
rect 253938 570480 253994 570489
rect 253938 570415 253994 570424
rect 253952 570042 253980 570415
rect 253940 570036 253992 570042
rect 253940 569978 253992 569984
rect 253388 569220 253440 569226
rect 253388 569162 253440 569168
rect 253296 565140 253348 565146
rect 253296 565082 253348 565088
rect 254596 563718 254624 652287
rect 257344 645924 257396 645930
rect 257344 645866 257396 645872
rect 254674 617264 254730 617273
rect 254674 617199 254730 617208
rect 254584 563712 254636 563718
rect 254584 563654 254636 563660
rect 254582 558784 254638 558793
rect 254582 558719 254638 558728
rect 254596 557598 254624 558719
rect 254584 557592 254636 557598
rect 254584 557534 254636 557540
rect 253204 555484 253256 555490
rect 253204 555426 253256 555432
rect 254398 552936 254454 552945
rect 254398 552871 254454 552880
rect 254412 551342 254440 552871
rect 254400 551336 254452 551342
rect 254400 551278 254452 551284
rect 254490 547088 254546 547097
rect 254490 547023 254546 547032
rect 254504 538214 254532 547023
rect 254688 541686 254716 617199
rect 254766 593872 254822 593881
rect 254766 593807 254822 593816
rect 254780 593434 254808 593807
rect 254768 593428 254820 593434
rect 254768 593370 254820 593376
rect 255964 581324 256016 581330
rect 255964 581266 256016 581272
rect 254676 541680 254728 541686
rect 254676 541622 254728 541628
rect 254582 541240 254638 541249
rect 254582 541175 254584 541184
rect 254636 541175 254638 541184
rect 254584 541146 254636 541152
rect 254504 538186 254624 538214
rect 254214 529544 254270 529553
rect 254214 529479 254270 529488
rect 254228 528630 254256 529479
rect 254216 528624 254268 528630
rect 254216 528566 254268 528572
rect 254030 523696 254086 523705
rect 254030 523631 254086 523640
rect 254044 523054 254072 523631
rect 254032 523048 254084 523054
rect 254032 522990 254084 522996
rect 254490 517848 254546 517857
rect 254490 517783 254546 517792
rect 254504 517546 254532 517783
rect 254492 517540 254544 517546
rect 254492 517482 254544 517488
rect 254398 512000 254454 512009
rect 254398 511935 254454 511944
rect 254412 510678 254440 511935
rect 254400 510672 254452 510678
rect 254400 510614 254452 510620
rect 254306 506152 254362 506161
rect 254306 506087 254362 506096
rect 254320 505170 254348 506087
rect 254308 505164 254360 505170
rect 254308 505106 254360 505112
rect 254214 500304 254270 500313
rect 254214 500239 254270 500248
rect 254228 499934 254256 500239
rect 254216 499928 254268 499934
rect 254216 499870 254268 499876
rect 254596 498846 254624 538186
rect 254674 535392 254730 535401
rect 254674 535327 254730 535336
rect 254688 534138 254716 535327
rect 254676 534132 254728 534138
rect 254676 534074 254728 534080
rect 254584 498840 254636 498846
rect 254584 498782 254636 498788
rect 254676 497548 254728 497554
rect 254676 497490 254728 497496
rect 254582 494456 254638 494465
rect 254582 494391 254638 494400
rect 254596 494086 254624 494391
rect 254584 494080 254636 494086
rect 254584 494022 254636 494028
rect 254688 489914 254716 497490
rect 254596 489886 254716 489914
rect 51724 485852 51776 485858
rect 51724 485794 51776 485800
rect 51354 397896 51410 397905
rect 51354 397831 51410 397840
rect 51354 356960 51410 356969
rect 51354 356895 51410 356904
rect 51368 282033 51396 356895
rect 51446 339416 51502 339425
rect 51446 339351 51502 339360
rect 51354 282024 51410 282033
rect 51354 281959 51410 281968
rect 51460 280809 51488 339351
rect 51630 333568 51686 333577
rect 51630 333503 51686 333512
rect 51538 310176 51594 310185
rect 51538 310111 51594 310120
rect 51552 281897 51580 310111
rect 51538 281888 51594 281897
rect 51538 281823 51594 281832
rect 51446 280800 51502 280809
rect 51446 280735 51502 280744
rect 51644 280673 51672 333503
rect 51630 280664 51686 280673
rect 51630 280599 51686 280608
rect 51736 201482 51764 485794
rect 254398 482760 254454 482769
rect 254398 482695 254454 482704
rect 254412 481710 254440 482695
rect 254400 481704 254452 481710
rect 254400 481646 254452 481652
rect 254214 476912 254270 476921
rect 254214 476847 254270 476856
rect 254228 476134 254256 476847
rect 254216 476128 254268 476134
rect 254216 476070 254268 476076
rect 254490 471064 254546 471073
rect 254490 470999 254546 471008
rect 254504 470626 254532 470999
rect 254492 470620 254544 470626
rect 254492 470562 254544 470568
rect 254306 459368 254362 459377
rect 254306 459303 254362 459312
rect 254320 458250 254348 459303
rect 254308 458244 254360 458250
rect 254308 458186 254360 458192
rect 254398 441824 254454 441833
rect 254398 441759 254400 441768
rect 254452 441759 254454 441768
rect 254400 441730 254452 441736
rect 254214 430128 254270 430137
rect 254214 430063 254270 430072
rect 254228 429214 254256 430063
rect 254216 429208 254268 429214
rect 254216 429150 254268 429156
rect 254398 418432 254454 418441
rect 254398 418367 254454 418376
rect 254412 418198 254440 418367
rect 254400 418192 254452 418198
rect 254400 418134 254452 418140
rect 254306 406736 254362 406745
rect 254306 406671 254362 406680
rect 254320 405754 254348 406671
rect 254308 405748 254360 405754
rect 254308 405690 254360 405696
rect 254490 400888 254546 400897
rect 254490 400823 254546 400832
rect 254504 400246 254532 400823
rect 254492 400240 254544 400246
rect 254492 400182 254544 400188
rect 254490 395040 254546 395049
rect 254490 394975 254492 394984
rect 254544 394975 254546 394984
rect 254492 394946 254544 394952
rect 254492 389224 254544 389230
rect 254490 389192 254492 389201
rect 254544 389192 254546 389201
rect 254490 389127 254546 389136
rect 254214 383344 254270 383353
rect 254214 383279 254270 383288
rect 254228 382294 254256 383279
rect 254216 382288 254268 382294
rect 254216 382230 254268 382236
rect 254122 377496 254178 377505
rect 254122 377431 254178 377440
rect 254136 376786 254164 377431
rect 254124 376780 254176 376786
rect 254124 376722 254176 376728
rect 254398 371648 254454 371657
rect 254398 371583 254454 371592
rect 254412 371278 254440 371583
rect 254400 371272 254452 371278
rect 254400 371214 254452 371220
rect 254490 365800 254546 365809
rect 254490 365735 254492 365744
rect 254544 365735 254546 365744
rect 254492 365706 254544 365712
rect 253938 359952 253994 359961
rect 253938 359887 253994 359896
rect 253952 358902 253980 359887
rect 253940 358896 253992 358902
rect 253940 358838 253992 358844
rect 254490 354104 254546 354113
rect 254490 354039 254546 354048
rect 254504 353326 254532 354039
rect 254492 353320 254544 353326
rect 254492 353262 254544 353268
rect 253386 332072 253442 332081
rect 253386 332007 253442 332016
rect 253202 331664 253258 331673
rect 253202 331599 253258 331608
rect 52090 286512 52146 286521
rect 52090 286447 52146 286456
rect 51908 281308 51960 281314
rect 51908 281250 51960 281256
rect 51920 280838 51948 281250
rect 52104 281246 52132 286447
rect 52920 281852 52972 281858
rect 52920 281794 52972 281800
rect 52092 281240 52144 281246
rect 52092 281182 52144 281188
rect 52932 281110 52960 281794
rect 54484 281308 54536 281314
rect 54484 281250 54536 281256
rect 55864 281308 55916 281314
rect 55864 281250 55916 281256
rect 52920 281104 52972 281110
rect 52920 281046 52972 281052
rect 51908 280832 51960 280838
rect 51908 280774 51960 280780
rect 53104 280832 53156 280838
rect 53104 280774 53156 280780
rect 52460 250504 52512 250510
rect 52460 250446 52512 250452
rect 51724 201476 51776 201482
rect 51724 201418 51776 201424
rect 51264 140752 51316 140758
rect 51264 140694 51316 140700
rect 52472 16574 52500 250446
rect 53116 157350 53144 280774
rect 53104 157344 53156 157350
rect 53104 157286 53156 157292
rect 54496 153202 54524 281250
rect 55876 280974 55904 281250
rect 55864 280968 55916 280974
rect 55864 280910 55916 280916
rect 59544 279472 59596 279478
rect 59544 279414 59596 279420
rect 54574 278760 54630 278769
rect 54574 278695 54630 278704
rect 54588 161430 54616 278695
rect 59358 278080 59414 278089
rect 59358 278015 59414 278024
rect 58992 262880 59044 262886
rect 58992 262822 59044 262828
rect 58900 261520 58952 261526
rect 58900 261462 58952 261468
rect 57060 233980 57112 233986
rect 57060 233922 57112 233928
rect 55862 223544 55918 223553
rect 55862 223479 55918 223488
rect 55876 164393 55904 223479
rect 57072 217433 57100 233922
rect 57428 228404 57480 228410
rect 57428 228346 57480 228352
rect 57336 222896 57388 222902
rect 57336 222838 57388 222844
rect 57244 221536 57296 221542
rect 57244 221478 57296 221484
rect 57152 220244 57204 220250
rect 57152 220186 57204 220192
rect 57058 217424 57114 217433
rect 57058 217359 57114 217368
rect 57164 209273 57192 220186
rect 57256 214606 57284 221478
rect 57244 214600 57296 214606
rect 57244 214542 57296 214548
rect 57150 209264 57206 209273
rect 57150 209199 57206 209208
rect 57348 205193 57376 222838
rect 57334 205184 57390 205193
rect 57334 205119 57390 205128
rect 57336 201476 57388 201482
rect 57336 201418 57388 201424
rect 57348 201113 57376 201418
rect 57334 201104 57390 201113
rect 57334 201039 57390 201048
rect 57336 197328 57388 197334
rect 57336 197270 57388 197276
rect 57348 197033 57376 197270
rect 57334 197024 57390 197033
rect 57334 196959 57390 196968
rect 57242 192944 57298 192953
rect 57242 192879 57298 192888
rect 57256 192506 57284 192879
rect 57244 192500 57296 192506
rect 57244 192442 57296 192448
rect 57336 189032 57388 189038
rect 57336 188974 57388 188980
rect 57348 188873 57376 188974
rect 57334 188864 57390 188873
rect 57334 188799 57390 188808
rect 56692 184884 56744 184890
rect 56692 184826 56744 184832
rect 56704 184793 56732 184826
rect 56690 184784 56746 184793
rect 56690 184719 56746 184728
rect 56692 180804 56744 180810
rect 56692 180746 56744 180752
rect 56704 180713 56732 180746
rect 56690 180704 56746 180713
rect 56690 180639 56746 180648
rect 57336 176656 57388 176662
rect 57334 176624 57336 176633
rect 57388 176624 57390 176633
rect 57334 176559 57390 176568
rect 57244 173392 57296 173398
rect 57244 173334 57296 173340
rect 57256 172553 57284 173334
rect 57242 172544 57298 172553
rect 57242 172479 57298 172488
rect 57336 169720 57388 169726
rect 57336 169662 57388 169668
rect 57348 168473 57376 169662
rect 57334 168464 57390 168473
rect 57334 168399 57390 168408
rect 55862 164384 55918 164393
rect 55862 164319 55918 164328
rect 54576 161424 54628 161430
rect 54576 161366 54628 161372
rect 57060 161424 57112 161430
rect 57060 161366 57112 161372
rect 57072 160313 57100 161366
rect 57058 160304 57114 160313
rect 57058 160239 57114 160248
rect 57060 157344 57112 157350
rect 57060 157286 57112 157292
rect 57072 156233 57100 157286
rect 57058 156224 57114 156233
rect 57058 156159 57114 156168
rect 54484 153196 54536 153202
rect 54484 153138 54536 153144
rect 57336 153196 57388 153202
rect 57336 153138 57388 153144
rect 57348 152153 57376 153138
rect 57334 152144 57390 152153
rect 57334 152079 57390 152088
rect 57336 149048 57388 149054
rect 57336 148990 57388 148996
rect 57348 148073 57376 148990
rect 57334 148064 57390 148073
rect 57334 147999 57390 148008
rect 57336 144560 57388 144566
rect 57336 144502 57388 144508
rect 57348 143993 57376 144502
rect 57334 143984 57390 143993
rect 57334 143919 57390 143928
rect 57440 142154 57468 228346
rect 57704 227044 57756 227050
rect 57704 226986 57756 226992
rect 57612 218748 57664 218754
rect 57612 218690 57664 218696
rect 57520 214600 57572 214606
rect 57520 214542 57572 214548
rect 57348 142126 57468 142154
rect 57348 135833 57376 142126
rect 57428 140752 57480 140758
rect 57428 140694 57480 140700
rect 57440 139913 57468 140694
rect 57426 139904 57482 139913
rect 57426 139839 57482 139848
rect 57334 135824 57390 135833
rect 57334 135759 57390 135768
rect 57532 123593 57560 214542
rect 57518 123584 57574 123593
rect 57518 123519 57574 123528
rect 57624 107273 57652 218690
rect 57610 107264 57666 107273
rect 57610 107199 57666 107208
rect 57716 103193 57744 226986
rect 58808 225752 58860 225758
rect 58808 225694 58860 225700
rect 57796 222964 57848 222970
rect 57796 222906 57848 222912
rect 57702 103184 57758 103193
rect 57702 103119 57758 103128
rect 57808 86873 57836 222906
rect 57888 218816 57940 218822
rect 57888 218758 57940 218764
rect 57794 86864 57850 86873
rect 57794 86799 57850 86808
rect 57900 78713 57928 218758
rect 58820 119513 58848 225694
rect 58912 127673 58940 261462
rect 58898 127664 58954 127673
rect 58898 127599 58954 127608
rect 58806 119504 58862 119513
rect 58806 119439 58862 119448
rect 59004 111353 59032 262822
rect 59268 260160 59320 260166
rect 59268 260102 59320 260108
rect 59084 236700 59136 236706
rect 59084 236642 59136 236648
rect 58990 111344 59046 111353
rect 58990 111279 59046 111288
rect 59096 82793 59124 236642
rect 59176 227112 59228 227118
rect 59176 227054 59228 227060
rect 59082 82784 59138 82793
rect 59082 82719 59138 82728
rect 57886 78704 57942 78713
rect 57886 78639 57942 78648
rect 59188 62393 59216 227054
rect 59280 90953 59308 260102
rect 59266 90944 59322 90953
rect 59266 90879 59322 90888
rect 59372 70553 59400 278015
rect 59450 276720 59506 276729
rect 59450 276655 59506 276664
rect 59464 95033 59492 276655
rect 59556 115433 59584 279414
rect 59728 232552 59780 232558
rect 59728 232494 59780 232500
rect 59636 229764 59688 229770
rect 59636 229706 59688 229712
rect 59542 115424 59598 115433
rect 59542 115359 59598 115368
rect 59450 95024 59506 95033
rect 59450 94959 59506 94968
rect 59358 70544 59414 70553
rect 59358 70479 59414 70488
rect 59648 66473 59676 229706
rect 59740 74633 59768 232494
rect 222844 222284 222896 222290
rect 222844 222226 222896 222232
rect 59820 221468 59872 221474
rect 59820 221410 59872 221416
rect 59832 99113 59860 221410
rect 60556 220176 60608 220182
rect 60556 220118 60608 220124
rect 60568 213897 60596 220118
rect 222856 215665 222884 222226
rect 224408 222216 224460 222222
rect 224408 222158 224460 222164
rect 222936 216708 222988 216714
rect 222936 216650 222988 216656
rect 222842 215656 222898 215665
rect 222842 215591 222898 215600
rect 60554 213888 60610 213897
rect 60554 213823 60610 213832
rect 222292 213036 222344 213042
rect 222292 212978 222344 212984
rect 222304 212809 222332 212978
rect 222290 212800 222346 212809
rect 222290 212735 222346 212744
rect 222948 207097 222976 216650
rect 223210 209944 223266 209953
rect 223210 209879 223266 209888
rect 222934 207088 222990 207097
rect 222934 207023 222990 207032
rect 223224 205630 223252 209879
rect 223212 205624 223264 205630
rect 223212 205566 223264 205572
rect 222842 204232 222898 204241
rect 222842 204167 222898 204176
rect 222856 190466 222884 204167
rect 223026 201376 223082 201385
rect 223026 201311 223082 201320
rect 222934 198520 222990 198529
rect 222934 198455 222990 198464
rect 222844 190460 222896 190466
rect 222844 190402 222896 190408
rect 222842 189952 222898 189961
rect 222842 189887 222898 189896
rect 222856 189106 222884 189887
rect 222844 189100 222896 189106
rect 222844 189042 222896 189048
rect 222842 187096 222898 187105
rect 222842 187031 222898 187040
rect 222856 186386 222884 187031
rect 222844 186380 222896 186386
rect 222844 186322 222896 186328
rect 222948 186318 222976 198455
rect 223040 189038 223068 201311
rect 224316 197396 224368 197402
rect 224316 197338 224368 197344
rect 224224 196036 224276 196042
rect 224224 195978 224276 195984
rect 223486 195664 223542 195673
rect 223486 195599 223542 195608
rect 223500 194614 223528 195599
rect 223488 194608 223540 194614
rect 223488 194550 223540 194556
rect 223486 192808 223542 192817
rect 223486 192743 223542 192752
rect 223500 191894 223528 192743
rect 223488 191888 223540 191894
rect 223488 191830 223540 191836
rect 223028 189032 223080 189038
rect 223028 188974 223080 188980
rect 222936 186312 222988 186318
rect 222936 186254 222988 186260
rect 222290 184240 222346 184249
rect 222290 184175 222346 184184
rect 222304 183802 222332 184175
rect 222292 183796 222344 183802
rect 222292 183738 222344 183744
rect 223486 181384 223542 181393
rect 223486 181319 223542 181328
rect 222658 178528 222714 178537
rect 222658 178463 222714 178472
rect 222672 176662 222700 178463
rect 223500 178022 223528 181319
rect 223488 178016 223540 178022
rect 223488 177958 223540 177964
rect 222660 176656 222712 176662
rect 222660 176598 222712 176604
rect 222658 175672 222714 175681
rect 222658 175607 222714 175616
rect 222672 175234 222700 175607
rect 222660 175228 222712 175234
rect 222660 175170 222712 175176
rect 222384 173188 222436 173194
rect 222384 173130 222436 173136
rect 222396 172825 222424 173130
rect 222382 172816 222438 172825
rect 222382 172751 222438 172760
rect 222476 171148 222528 171154
rect 222476 171090 222528 171096
rect 222488 169969 222516 171090
rect 222474 169960 222530 169969
rect 222474 169895 222530 169904
rect 222936 169788 222988 169794
rect 222936 169730 222988 169736
rect 222948 167113 222976 169730
rect 222934 167104 222990 167113
rect 222934 167039 222990 167048
rect 223488 167068 223540 167074
rect 223488 167010 223540 167016
rect 223028 165640 223080 165646
rect 223028 165582 223080 165588
rect 222936 164280 222988 164286
rect 222936 164222 222988 164228
rect 222948 158545 222976 164222
rect 223040 161401 223068 165582
rect 223500 164257 223528 167010
rect 223486 164248 223542 164257
rect 223486 164183 223542 164192
rect 223488 162920 223540 162926
rect 223488 162862 223540 162868
rect 223026 161392 223082 161401
rect 223026 161327 223082 161336
rect 222934 158536 222990 158545
rect 222934 158471 222990 158480
rect 222568 157140 222620 157146
rect 222568 157082 222620 157088
rect 222580 152833 222608 157082
rect 223500 155689 223528 162862
rect 223486 155680 223542 155689
rect 223486 155615 223542 155624
rect 222936 154624 222988 154630
rect 222936 154566 222988 154572
rect 222844 153264 222896 153270
rect 222844 153206 222896 153212
rect 222566 152824 222622 152833
rect 222566 152759 222622 152768
rect 222476 144356 222528 144362
rect 222476 144298 222528 144304
rect 222488 144265 222516 144298
rect 222474 144256 222530 144265
rect 222474 144191 222530 144200
rect 222476 137284 222528 137290
rect 222476 137226 222528 137232
rect 222488 132841 222516 137226
rect 222856 135697 222884 153206
rect 222948 138553 222976 154566
rect 223488 150476 223540 150482
rect 223488 150418 223540 150424
rect 223500 149977 223528 150418
rect 223486 149968 223542 149977
rect 223486 149903 223542 149912
rect 223488 147280 223540 147286
rect 223488 147222 223540 147228
rect 223500 147121 223528 147222
rect 223486 147112 223542 147121
rect 223486 147047 223542 147056
rect 223488 141500 223540 141506
rect 223488 141442 223540 141448
rect 223500 141409 223528 141442
rect 223486 141400 223542 141409
rect 223486 141335 223542 141344
rect 222934 138544 222990 138553
rect 222934 138479 222990 138488
rect 222842 135688 222898 135697
rect 222842 135623 222898 135632
rect 223120 133204 223172 133210
rect 223120 133146 223172 133152
rect 222474 132832 222530 132841
rect 222474 132767 222530 132776
rect 223132 129985 223160 133146
rect 223488 130416 223540 130422
rect 223488 130358 223540 130364
rect 223118 129976 223174 129985
rect 223118 129911 223174 129920
rect 222476 128308 222528 128314
rect 222476 128250 222528 128256
rect 222488 124273 222516 128250
rect 223500 127129 223528 130358
rect 223486 127120 223542 127129
rect 223486 127055 223542 127064
rect 223212 124636 223264 124642
rect 223212 124578 223264 124584
rect 222474 124264 222530 124273
rect 222474 124199 222530 124208
rect 223224 121417 223252 124578
rect 223210 121408 223266 121417
rect 223210 121343 223266 121352
rect 223488 118652 223540 118658
rect 223488 118594 223540 118600
rect 223500 118561 223528 118594
rect 223486 118552 223542 118561
rect 223486 118487 223542 118496
rect 223488 115932 223540 115938
rect 223488 115874 223540 115880
rect 223500 115705 223528 115874
rect 223486 115696 223542 115705
rect 223486 115631 223542 115640
rect 222200 113008 222252 113014
rect 222200 112950 222252 112956
rect 222212 112849 222240 112950
rect 222198 112840 222254 112849
rect 222198 112775 222254 112784
rect 223488 110424 223540 110430
rect 223488 110366 223540 110372
rect 223500 109993 223528 110366
rect 223486 109984 223542 109993
rect 223486 109919 223542 109928
rect 222660 107636 222712 107642
rect 222660 107578 222712 107584
rect 222672 107137 222700 107578
rect 222658 107128 222714 107137
rect 222658 107063 222714 107072
rect 222844 104848 222896 104854
rect 222844 104790 222896 104796
rect 222856 104281 222884 104790
rect 222842 104272 222898 104281
rect 222842 104207 222898 104216
rect 223488 102128 223540 102134
rect 223488 102070 223540 102076
rect 223500 101425 223528 102070
rect 223486 101416 223542 101425
rect 223486 101351 223542 101360
rect 223028 99340 223080 99346
rect 223028 99282 223080 99288
rect 59818 99104 59874 99113
rect 59818 99039 59874 99048
rect 223040 98569 223068 99282
rect 223026 98560 223082 98569
rect 223026 98495 223082 98504
rect 223120 96620 223172 96626
rect 223120 96562 223172 96568
rect 223132 95713 223160 96562
rect 223118 95704 223174 95713
rect 223118 95639 223174 95648
rect 223488 93832 223540 93838
rect 223488 93774 223540 93780
rect 223500 92857 223528 93774
rect 223486 92848 223542 92857
rect 223486 92783 223542 92792
rect 223396 91792 223448 91798
rect 223396 91734 223448 91740
rect 223408 87145 223436 91734
rect 223488 90364 223540 90370
rect 223488 90306 223540 90312
rect 223500 90001 223528 90306
rect 223486 89992 223542 90001
rect 223486 89927 223542 89936
rect 223488 87644 223540 87650
rect 223488 87586 223540 87592
rect 223394 87136 223450 87145
rect 223394 87071 223450 87080
rect 223500 84289 223528 87586
rect 223486 84280 223542 84289
rect 223486 84215 223542 84224
rect 223486 81424 223542 81433
rect 223486 81359 223488 81368
rect 223540 81359 223542 81368
rect 223488 81330 223540 81336
rect 222476 78600 222528 78606
rect 222474 78568 222476 78577
rect 222528 78568 222530 78577
rect 222474 78503 222530 78512
rect 222200 75744 222252 75750
rect 222198 75712 222200 75721
rect 222252 75712 222254 75721
rect 222198 75647 222254 75656
rect 59726 74624 59782 74633
rect 59726 74559 59782 74568
rect 224236 73098 224264 195978
rect 224328 75750 224356 197338
rect 224420 113014 224448 222158
rect 226064 220856 226116 220862
rect 226064 220798 226116 220804
rect 226076 213042 226104 220798
rect 253216 218822 253244 331599
rect 253400 221542 253428 332007
rect 253570 331392 253626 331401
rect 253570 331327 253626 331336
rect 253584 222970 253612 331327
rect 254214 330712 254270 330721
rect 254214 330647 254270 330656
rect 254228 329934 254256 330647
rect 254216 329928 254268 329934
rect 254216 329870 254268 329876
rect 254492 325644 254544 325650
rect 254492 325586 254544 325592
rect 254504 324873 254532 325586
rect 254490 324864 254546 324873
rect 254490 324799 254546 324808
rect 254308 320136 254360 320142
rect 254308 320078 254360 320084
rect 254320 319025 254348 320078
rect 254306 319016 254362 319025
rect 254306 318951 254362 318960
rect 254214 307320 254270 307329
rect 254214 307255 254270 307264
rect 254228 306406 254256 307255
rect 254216 306400 254268 306406
rect 254216 306342 254268 306348
rect 254030 289776 254086 289785
rect 254030 289711 254086 289720
rect 254044 280974 254072 289711
rect 254306 283928 254362 283937
rect 254306 283863 254362 283872
rect 254320 282946 254348 283863
rect 254308 282940 254360 282946
rect 254308 282882 254360 282888
rect 254032 280968 254084 280974
rect 254032 280910 254084 280916
rect 253572 222964 253624 222970
rect 253572 222906 253624 222912
rect 254596 222902 254624 489886
rect 254674 488608 254730 488617
rect 254674 488543 254676 488552
rect 254728 488543 254730 488552
rect 254676 488514 254728 488520
rect 254674 465216 254730 465225
rect 254674 465151 254730 465160
rect 254688 465118 254716 465151
rect 254676 465112 254728 465118
rect 254676 465054 254728 465060
rect 254674 453520 254730 453529
rect 254674 453455 254730 453464
rect 254688 452674 254716 453455
rect 254676 452668 254728 452674
rect 254676 452610 254728 452616
rect 254674 447672 254730 447681
rect 254674 447607 254730 447616
rect 254688 447166 254716 447607
rect 254676 447160 254728 447166
rect 254676 447102 254728 447108
rect 254674 435976 254730 435985
rect 254674 435911 254730 435920
rect 254688 434790 254716 435911
rect 254676 434784 254728 434790
rect 254676 434726 254728 434732
rect 254674 424280 254730 424289
rect 254674 424215 254730 424224
rect 254688 423706 254716 424215
rect 254676 423700 254728 423706
rect 254676 423642 254728 423648
rect 254674 412584 254730 412593
rect 254674 412519 254730 412528
rect 254688 345014 254716 412519
rect 254766 348256 254822 348265
rect 254766 348191 254822 348200
rect 254780 347818 254808 348191
rect 254768 347812 254820 347818
rect 254768 347754 254820 347760
rect 254688 344986 254808 345014
rect 254674 342408 254730 342417
rect 254674 342343 254730 342352
rect 254688 342310 254716 342343
rect 254676 342304 254728 342310
rect 254676 342246 254728 342252
rect 254674 336560 254730 336569
rect 254674 336495 254730 336504
rect 254688 335374 254716 336495
rect 254780 336054 254808 344986
rect 254768 336048 254820 336054
rect 254768 335990 254820 335996
rect 254676 335368 254728 335374
rect 254676 335310 254728 335316
rect 254676 329860 254728 329866
rect 254676 329802 254728 329808
rect 254688 313177 254716 329802
rect 254674 313168 254730 313177
rect 254674 313103 254730 313112
rect 254674 301472 254730 301481
rect 254674 301407 254730 301416
rect 254688 300898 254716 301407
rect 254676 300892 254728 300898
rect 254676 300834 254728 300840
rect 254674 295624 254730 295633
rect 254674 295559 254730 295568
rect 254688 295390 254716 295559
rect 254676 295384 254728 295390
rect 254676 295326 254728 295332
rect 254584 222896 254636 222902
rect 254584 222838 254636 222844
rect 253388 221536 253440 221542
rect 253388 221478 253440 221484
rect 253204 218816 253256 218822
rect 253204 218758 253256 218764
rect 247684 215348 247736 215354
rect 247684 215290 247736 215296
rect 246304 213988 246356 213994
rect 246304 213930 246356 213936
rect 226064 213036 226116 213042
rect 226064 212978 226116 212984
rect 243544 212560 243596 212566
rect 243544 212502 243596 212508
rect 242164 211200 242216 211206
rect 242164 211142 242216 211148
rect 239404 209840 239456 209846
rect 239404 209782 239456 209788
rect 238024 208412 238076 208418
rect 238024 208354 238076 208360
rect 232504 207052 232556 207058
rect 232504 206994 232556 207000
rect 229744 205692 229796 205698
rect 229744 205634 229796 205640
rect 228364 200184 228416 200190
rect 228364 200126 228416 200132
rect 225604 198756 225656 198762
rect 225604 198698 225656 198704
rect 224960 189100 225012 189106
rect 224960 189042 225012 189048
rect 224972 182170 225000 189042
rect 224960 182164 225012 182170
rect 224960 182106 225012 182112
rect 224408 113008 224460 113014
rect 224408 112950 224460 112956
rect 225616 78606 225644 198698
rect 225788 183796 225840 183802
rect 225788 183738 225840 183744
rect 225800 179382 225828 183738
rect 225788 179376 225840 179382
rect 225788 179318 225840 179324
rect 225696 157412 225748 157418
rect 225696 157354 225748 157360
rect 225708 144362 225736 157354
rect 225696 144356 225748 144362
rect 225696 144298 225748 144304
rect 228376 81394 228404 200126
rect 228456 186380 228508 186386
rect 228456 186322 228508 186328
rect 228468 180810 228496 186322
rect 228456 180804 228508 180810
rect 228456 180746 228508 180752
rect 229100 161492 229152 161498
rect 229100 161434 229152 161440
rect 228456 158772 228508 158778
rect 228456 158714 228508 158720
rect 228468 147286 228496 158714
rect 229112 157146 229140 161434
rect 229100 157140 229152 157146
rect 229100 157082 229152 157088
rect 228456 147280 228508 147286
rect 228456 147222 228508 147228
rect 228456 144968 228508 144974
rect 228456 144910 228508 144916
rect 228468 124642 228496 144910
rect 228456 124636 228508 124642
rect 228456 124578 228508 124584
rect 229756 90370 229784 205634
rect 229836 205624 229888 205630
rect 229836 205566 229888 205572
rect 229848 193186 229876 205566
rect 229836 193180 229888 193186
rect 229836 193122 229888 193128
rect 229928 191888 229980 191894
rect 229928 191830 229980 191836
rect 229940 183530 229968 191830
rect 229928 183524 229980 183530
rect 229928 183466 229980 183472
rect 231124 160132 231176 160138
rect 231124 160074 231176 160080
rect 229836 155984 229888 155990
rect 229836 155926 229888 155932
rect 229848 141506 229876 155926
rect 231136 150482 231164 160074
rect 231124 150476 231176 150482
rect 231124 150418 231176 150424
rect 231124 146328 231176 146334
rect 231124 146270 231176 146276
rect 229836 141500 229888 141506
rect 229836 141442 229888 141448
rect 231136 128314 231164 146270
rect 231124 128308 231176 128314
rect 231124 128250 231176 128256
rect 232516 93838 232544 206994
rect 233976 194608 234028 194614
rect 233976 194550 234028 194556
rect 233884 190528 233936 190534
rect 233884 190470 233936 190476
rect 232596 143608 232648 143614
rect 232596 143550 232648 143556
rect 232608 118658 232636 143550
rect 232596 118652 232648 118658
rect 232596 118594 232648 118600
rect 232504 93832 232556 93838
rect 232504 93774 232556 93780
rect 229744 90364 229796 90370
rect 229744 90306 229796 90312
rect 228364 81388 228416 81394
rect 228364 81330 228416 81336
rect 225604 78600 225656 78606
rect 225604 78542 225656 78548
rect 224316 75744 224368 75750
rect 224316 75686 224368 75692
rect 222200 73092 222252 73098
rect 222200 73034 222252 73040
rect 224224 73092 224276 73098
rect 224224 73034 224276 73040
rect 222212 72865 222240 73034
rect 222198 72856 222254 72865
rect 222198 72791 222254 72800
rect 223488 70372 223540 70378
rect 223488 70314 223540 70320
rect 223500 70009 223528 70314
rect 223486 70000 223542 70009
rect 223486 69935 223542 69944
rect 223488 67584 223540 67590
rect 223488 67526 223540 67532
rect 223500 67153 223528 67526
rect 223486 67144 223542 67153
rect 223486 67079 223542 67088
rect 59634 66464 59690 66473
rect 59634 66399 59690 66408
rect 233896 64870 233924 190470
rect 233988 184890 234016 194550
rect 235264 193248 235316 193254
rect 235264 193190 235316 193196
rect 233976 184884 234028 184890
rect 233976 184826 234028 184832
rect 233976 147688 234028 147694
rect 233976 147630 234028 147636
rect 233988 130422 234016 147630
rect 233976 130416 234028 130422
rect 233976 130358 234028 130364
rect 235276 67590 235304 193190
rect 236644 151836 236696 151842
rect 236644 151778 236696 151784
rect 235356 149116 235408 149122
rect 235356 149058 235408 149064
rect 235368 133210 235396 149058
rect 236656 137290 236684 151778
rect 236644 137284 236696 137290
rect 236644 137226 236696 137232
rect 235356 133204 235408 133210
rect 235356 133146 235408 133152
rect 238036 96626 238064 208354
rect 239416 99346 239444 209782
rect 242176 102134 242204 211142
rect 243556 104854 243584 212502
rect 246316 107642 246344 213930
rect 247696 110430 247724 215290
rect 250444 194608 250496 194614
rect 250444 194550 250496 194556
rect 247684 110424 247736 110430
rect 247684 110366 247736 110372
rect 246304 107636 246356 107642
rect 246304 107578 246356 107584
rect 243544 104848 243596 104854
rect 243544 104790 243596 104796
rect 242164 102128 242216 102134
rect 242164 102070 242216 102076
rect 239404 99340 239456 99346
rect 239404 99282 239456 99288
rect 238024 96620 238076 96626
rect 238024 96562 238076 96568
rect 250456 70378 250484 194550
rect 251824 142180 251876 142186
rect 251824 142122 251876 142128
rect 251836 115938 251864 142122
rect 251824 115932 251876 115938
rect 251824 115874 251876 115880
rect 255976 75886 256004 581266
rect 256056 570036 256108 570042
rect 256056 569978 256108 569984
rect 255964 75880 256016 75886
rect 255964 75822 256016 75828
rect 256068 73166 256096 569978
rect 256148 358896 256200 358902
rect 256148 358838 256200 358844
rect 256160 306338 256188 358838
rect 256148 306332 256200 306338
rect 256148 306274 256200 306280
rect 257356 142118 257384 645866
rect 257448 543046 257476 660554
rect 264244 622464 264296 622470
rect 264244 622406 264296 622412
rect 260104 587988 260156 587994
rect 260104 587930 260156 587936
rect 257436 543040 257488 543046
rect 257436 542982 257488 542988
rect 257436 499928 257488 499934
rect 257436 499870 257488 499876
rect 257344 142112 257396 142118
rect 257344 142054 257396 142060
rect 257448 128314 257476 499870
rect 258724 497752 258776 497758
rect 258724 497694 258776 497700
rect 257620 497616 257672 497622
rect 257620 497558 257672 497564
rect 257528 441788 257580 441794
rect 257528 441730 257580 441736
rect 257436 128308 257488 128314
rect 257436 128250 257488 128256
rect 257540 113150 257568 441730
rect 257632 218657 257660 497558
rect 258080 349852 258132 349858
rect 258080 349794 258132 349800
rect 257618 218648 257674 218657
rect 257618 218583 257674 218592
rect 257528 113144 257580 113150
rect 257528 113086 257580 113092
rect 256056 73160 256108 73166
rect 256056 73102 256108 73108
rect 250444 70372 250496 70378
rect 250444 70314 250496 70320
rect 235264 67584 235316 67590
rect 235264 67526 235316 67532
rect 222844 64864 222896 64870
rect 222844 64806 222896 64812
rect 233884 64864 233936 64870
rect 233884 64806 233936 64812
rect 222856 64297 222884 64806
rect 222842 64288 222898 64297
rect 222842 64223 222898 64232
rect 59174 62384 59230 62393
rect 59174 62319 59230 62328
rect 215300 61600 215352 61606
rect 215300 61542 215352 61548
rect 168380 61532 168432 61538
rect 168380 61474 168432 61480
rect 158720 61464 158772 61470
rect 126978 61432 127034 61441
rect 158720 61406 158772 61412
rect 126978 61367 127034 61376
rect 154580 61396 154632 61402
rect 99380 43444 99432 43450
rect 99380 43386 99432 43392
rect 56600 40724 56652 40730
rect 56600 40666 56652 40672
rect 56612 16574 56640 40666
rect 70400 33788 70452 33794
rect 70400 33730 70452 33736
rect 60740 21412 60792 21418
rect 60740 21354 60792 21360
rect 60752 16574 60780 21354
rect 70412 16574 70440 33730
rect 77300 29640 77352 29646
rect 77300 29582 77352 29588
rect 77312 16574 77340 29582
rect 92480 26920 92532 26926
rect 92480 26862 92532 26868
rect 52472 16546 53328 16574
rect 56612 16546 56824 16574
rect 60752 16546 60872 16574
rect 70412 16546 71544 16574
rect 77312 16546 78168 16574
rect 46664 6316 46716 6322
rect 46664 6258 46716 6264
rect 46676 480 46704 6258
rect 50160 4888 50212 4894
rect 50160 4830 50212 4836
rect 50172 480 50200 4830
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 60844 480 60872 16546
rect 67916 7744 67968 7750
rect 67916 7686 67968 7692
rect 64328 7676 64380 7682
rect 64328 7618 64380 7624
rect 64340 480 64368 7618
rect 67928 480 67956 7686
rect 71516 480 71544 16546
rect 74998 8936 75054 8945
rect 74998 8871 75054 8880
rect 75012 480 75040 8871
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 81624 15904 81676 15910
rect 81624 15846 81676 15852
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 15846
rect 89168 9036 89220 9042
rect 89168 8978 89220 8984
rect 85672 8968 85724 8974
rect 85672 8910 85724 8916
rect 85684 480 85712 8910
rect 89180 480 89208 8978
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 26862
rect 99392 16574 99420 43386
rect 120080 40792 120132 40798
rect 120080 40734 120132 40740
rect 113180 37936 113232 37942
rect 113180 37878 113232 37884
rect 110420 35284 110472 35290
rect 110420 35226 110472 35232
rect 102140 19984 102192 19990
rect 102140 19926 102192 19932
rect 99392 16546 99880 16574
rect 95790 10296 95846 10305
rect 95790 10231 95846 10240
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 95804 354 95832 10231
rect 99852 480 99880 16546
rect 102152 3602 102180 19926
rect 106280 18692 106332 18698
rect 106280 18634 106332 18640
rect 106292 16574 106320 18634
rect 110432 16574 110460 35226
rect 113192 16574 113220 37878
rect 117320 36576 117372 36582
rect 117320 36518 117372 36524
rect 106292 16546 106504 16574
rect 110432 16546 110552 16574
rect 113192 16546 114048 16574
rect 102140 3596 102192 3602
rect 102140 3538 102192 3544
rect 103336 3596 103388 3602
rect 103336 3538 103388 3544
rect 103348 480 103376 3538
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 110524 480 110552 16546
rect 114020 480 114048 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117332 354 117360 36518
rect 120092 16574 120120 40734
rect 120092 16546 120672 16574
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 124680 3596 124732 3602
rect 124680 3538 124732 3544
rect 124692 480 124720 3538
rect 126992 480 127020 61367
rect 154580 61338 154632 61344
rect 136638 60072 136694 60081
rect 136638 60007 136694 60016
rect 129738 59936 129794 59945
rect 129738 59871 129794 59880
rect 129752 16574 129780 59871
rect 133880 58676 133932 58682
rect 133880 58618 133932 58624
rect 129752 16546 130608 16574
rect 130580 480 130608 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 58618
rect 136652 16574 136680 60007
rect 147678 58576 147734 58585
rect 147678 58511 147734 58520
rect 147692 16574 147720 58511
rect 151820 42084 151872 42090
rect 151820 42026 151872 42032
rect 136652 16546 137232 16574
rect 147692 16546 147904 16574
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 143538 10432 143594 10441
rect 143538 10367 143594 10376
rect 141240 5024 141292 5030
rect 141240 4966 141292 4972
rect 141252 480 141280 4966
rect 143552 3398 143580 10367
rect 143540 3392 143592 3398
rect 143540 3334 143592 3340
rect 144736 3392 144788 3398
rect 144736 3334 144788 3340
rect 144748 480 144776 3334
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 151832 480 151860 42026
rect 154592 16574 154620 61338
rect 158732 16574 158760 61406
rect 165618 60208 165674 60217
rect 165618 60143 165674 60152
rect 165632 16574 165660 60143
rect 154592 16546 155448 16574
rect 158732 16546 158944 16574
rect 165632 16546 166120 16574
rect 155420 480 155448 16546
rect 158916 480 158944 16546
rect 162490 3360 162546 3369
rect 162490 3295 162546 3304
rect 162504 480 162532 3295
rect 166092 480 166120 16546
rect 168392 3398 168420 61474
rect 211160 60104 211212 60110
rect 211160 60046 211212 60052
rect 193220 60036 193272 60042
rect 193220 59978 193272 59984
rect 172520 58744 172572 58750
rect 172520 58686 172572 58692
rect 172532 16574 172560 58686
rect 190460 57316 190512 57322
rect 190460 57258 190512 57264
rect 176660 57248 176712 57254
rect 176660 57190 176712 57196
rect 172532 16546 172744 16574
rect 168380 3392 168432 3398
rect 168380 3334 168432 3340
rect 169576 3392 169628 3398
rect 169576 3334 169628 3340
rect 169588 480 169616 3334
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 176672 480 176700 57190
rect 179420 55888 179472 55894
rect 179420 55830 179472 55836
rect 179432 16574 179460 55830
rect 179432 16546 180288 16574
rect 180260 480 180288 16546
rect 187330 4856 187386 4865
rect 187330 4791 187386 4800
rect 183742 3496 183798 3505
rect 183742 3431 183798 3440
rect 183756 480 183784 3431
rect 187344 480 187372 4791
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173134 -960 173246 326
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 57258
rect 193232 3398 193260 59978
rect 204260 54528 204312 54534
rect 204260 54470 204312 54476
rect 201500 47592 201552 47598
rect 201500 47534 201552 47540
rect 197360 18760 197412 18766
rect 197360 18702 197412 18708
rect 197372 16574 197400 18702
rect 197372 16546 197952 16574
rect 193220 3392 193272 3398
rect 193220 3334 193272 3340
rect 194416 3392 194468 3398
rect 194416 3334 194468 3340
rect 194428 480 194456 3334
rect 197924 480 197952 16546
rect 201512 480 201540 47534
rect 204272 16574 204300 54470
rect 208400 40860 208452 40866
rect 208400 40802 208452 40808
rect 208412 16574 208440 40802
rect 211172 16574 211200 60046
rect 204272 16546 205128 16574
rect 208412 16546 208624 16574
rect 211172 16546 211752 16574
rect 205100 480 205128 16546
rect 208596 480 208624 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 61542
rect 229100 57384 229152 57390
rect 229100 57326 229152 57332
rect 226340 55956 226392 55962
rect 226340 55898 226392 55904
rect 218060 54596 218112 54602
rect 218060 54538 218112 54544
rect 218072 3398 218100 54538
rect 222752 3664 222804 3670
rect 222752 3606 222804 3612
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 219256 3392 219308 3398
rect 219256 3334 219308 3340
rect 219268 480 219296 3334
rect 222764 480 222792 3606
rect 226352 480 226380 55898
rect 229112 16574 229140 57326
rect 233240 56024 233292 56030
rect 233240 55966 233292 55972
rect 233252 16574 233280 55966
rect 247040 54664 247092 54670
rect 247040 54606 247092 54612
rect 236000 35352 236052 35358
rect 236000 35294 236052 35300
rect 236012 16574 236040 35294
rect 247052 16574 247080 54606
rect 251180 50380 251232 50386
rect 251180 50322 251232 50328
rect 229112 16546 229416 16574
rect 233252 16546 233464 16574
rect 236012 16546 236592 16574
rect 247052 16546 247632 16574
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 16546
rect 233436 480 233464 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 242900 10396 242952 10402
rect 242900 10338 242952 10344
rect 240140 10328 240192 10334
rect 240140 10270 240192 10276
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 354 240180 10270
rect 242912 3398 242940 10338
rect 242900 3392 242952 3398
rect 242900 3334 242952 3340
rect 244096 3392 244148 3398
rect 244096 3334 244148 3340
rect 244108 480 244136 3334
rect 247604 480 247632 16546
rect 251192 480 251220 50322
rect 258092 16574 258120 349794
rect 258736 228410 258764 497694
rect 258724 228404 258776 228410
rect 258724 228346 258776 228352
rect 260116 77246 260144 587930
rect 261484 575544 261536 575550
rect 261484 575486 261536 575492
rect 260196 541204 260248 541210
rect 260196 541146 260248 541152
rect 260208 89010 260236 541146
rect 260288 497684 260340 497690
rect 260288 497626 260340 497632
rect 260300 233986 260328 497626
rect 260380 395004 260432 395010
rect 260380 394946 260432 394952
rect 260392 307766 260420 394946
rect 260840 337408 260892 337414
rect 260840 337350 260892 337356
rect 260380 307760 260432 307766
rect 260380 307702 260432 307708
rect 260288 233980 260340 233986
rect 260288 233922 260340 233928
rect 260196 89004 260248 89010
rect 260196 88946 260248 88952
rect 260104 77240 260156 77246
rect 260104 77182 260156 77188
rect 260852 16574 260880 337350
rect 261496 74526 261524 575486
rect 261576 494080 261628 494086
rect 261576 494022 261628 494028
rect 261588 126954 261616 494022
rect 261576 126948 261628 126954
rect 261576 126890 261628 126896
rect 264256 90370 264284 622406
rect 264348 558210 264376 700470
rect 265624 700460 265676 700466
rect 265624 700402 265676 700408
rect 265636 559570 265664 700402
rect 267660 697678 267688 703520
rect 283852 700534 283880 703520
rect 283840 700528 283892 700534
rect 283840 700470 283892 700476
rect 300136 700466 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300124 700460 300176 700466
rect 300124 700402 300176 700408
rect 320916 700460 320968 700466
rect 320916 700402 320968 700408
rect 317420 700392 317472 700398
rect 317420 700334 317472 700340
rect 266360 697672 266412 697678
rect 266360 697614 266412 697620
rect 267648 697672 267700 697678
rect 267648 697614 267700 697620
rect 266372 592686 266400 697614
rect 316132 683188 316184 683194
rect 316132 683130 316184 683136
rect 279424 663128 279476 663134
rect 279424 663070 279476 663076
rect 279332 661768 279384 661774
rect 279332 661710 279384 661716
rect 278136 660544 278188 660550
rect 278136 660486 278188 660492
rect 273996 640348 274048 640354
rect 273996 640290 274048 640296
rect 271236 633480 271288 633486
rect 271236 633422 271288 633428
rect 269764 611380 269816 611386
rect 269764 611322 269816 611328
rect 266360 592680 266412 592686
rect 266360 592622 266412 592628
rect 265624 559564 265676 559570
rect 265624 559506 265676 559512
rect 264336 558204 264388 558210
rect 264336 558146 264388 558152
rect 265624 557592 265676 557598
rect 265624 557534 265676 557540
rect 264980 496120 265032 496126
rect 264980 496062 265032 496068
rect 264336 470620 264388 470626
rect 264336 470562 264388 470568
rect 264348 121446 264376 470562
rect 264428 282940 264480 282946
rect 264428 282882 264480 282888
rect 264336 121440 264388 121446
rect 264336 121382 264388 121388
rect 264244 90364 264296 90370
rect 264244 90306 264296 90312
rect 261484 74520 261536 74526
rect 261484 74462 261536 74468
rect 264440 62082 264468 282882
rect 264428 62076 264480 62082
rect 264428 62018 264480 62024
rect 258092 16546 258304 16574
rect 260852 16546 261800 16574
rect 254216 14476 254268 14482
rect 254216 14418 254268 14424
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 14418
rect 258276 480 258304 16546
rect 261772 480 261800 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 496062
rect 265636 70378 265664 557534
rect 268384 551336 268436 551342
rect 268384 551278 268436 551284
rect 267004 541680 267056 541686
rect 267004 541622 267056 541628
rect 265716 476128 265768 476134
rect 265716 476070 265768 476076
rect 265728 122806 265756 476070
rect 265716 122800 265768 122806
rect 265716 122742 265768 122748
rect 267016 85542 267044 541622
rect 267740 338836 267792 338842
rect 267740 338778 267792 338784
rect 267004 85536 267056 85542
rect 267004 85478 267056 85484
rect 265624 70372 265676 70378
rect 265624 70314 265676 70320
rect 267752 16574 267780 338778
rect 268396 69018 268424 551278
rect 268476 481704 268528 481710
rect 268476 481646 268528 481652
rect 268488 124166 268516 481646
rect 268476 124160 268528 124166
rect 268476 124102 268528 124108
rect 269776 84182 269804 611322
rect 271144 593428 271196 593434
rect 271144 593370 271196 593376
rect 269856 528624 269908 528630
rect 269856 528566 269908 528572
rect 269868 136610 269896 528566
rect 269948 458244 270000 458250
rect 269948 458186 270000 458192
rect 269856 136604 269908 136610
rect 269856 136546 269908 136552
rect 269960 118658 269988 458186
rect 269948 118652 270000 118658
rect 269948 118594 270000 118600
rect 269764 84176 269816 84182
rect 269764 84118 269816 84124
rect 271156 78674 271184 593370
rect 271248 139398 271276 633422
rect 273904 599004 273956 599010
rect 273904 598946 273956 598952
rect 271328 510672 271380 510678
rect 271328 510614 271380 510620
rect 271236 139392 271288 139398
rect 271236 139334 271288 139340
rect 271340 131102 271368 510614
rect 271880 344344 271932 344350
rect 271880 344286 271932 344292
rect 271328 131096 271380 131102
rect 271328 131038 271380 131044
rect 271144 78668 271196 78674
rect 271144 78610 271196 78616
rect 268384 69012 268436 69018
rect 268384 68954 268436 68960
rect 271892 16574 271920 344286
rect 273916 80034 273944 598946
rect 274008 140758 274036 640290
rect 278044 627972 278096 627978
rect 278044 627914 278096 627920
rect 275284 604512 275336 604518
rect 275284 604454 275336 604460
rect 274088 517540 274140 517546
rect 274088 517482 274140 517488
rect 273996 140752 274048 140758
rect 273996 140694 274048 140700
rect 274100 132462 274128 517482
rect 274088 132456 274140 132462
rect 274088 132398 274140 132404
rect 275296 82822 275324 604454
rect 276664 539640 276716 539646
rect 276664 539582 276716 539588
rect 275376 523048 275428 523054
rect 275376 522990 275428 522996
rect 275388 135250 275416 522990
rect 275468 505164 275520 505170
rect 275468 505106 275520 505112
rect 275376 135244 275428 135250
rect 275376 135186 275428 135192
rect 275480 129742 275508 505106
rect 276020 487824 276072 487830
rect 276020 487766 276072 487772
rect 275468 129736 275520 129742
rect 275468 129678 275520 129684
rect 275284 82816 275336 82822
rect 275284 82758 275336 82764
rect 273904 80028 273956 80034
rect 273904 79970 273956 79976
rect 267752 16546 268424 16574
rect 271892 16546 272472 16574
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 272444 480 272472 16546
rect 276032 480 276060 487766
rect 276676 281042 276704 539582
rect 276664 281036 276716 281042
rect 276664 280978 276716 280984
rect 278056 137970 278084 627914
rect 278148 543114 278176 660486
rect 279056 660272 279108 660278
rect 279056 660214 279108 660220
rect 278964 660136 279016 660142
rect 278964 660078 279016 660084
rect 278688 641164 278740 641170
rect 278688 641106 278740 641112
rect 278596 641028 278648 641034
rect 278596 640970 278648 640976
rect 278608 630057 278636 640970
rect 278594 630048 278650 630057
rect 278594 629983 278650 629992
rect 278700 610065 278728 641106
rect 278686 610056 278742 610065
rect 278686 609991 278742 610000
rect 278976 543658 279004 660078
rect 278964 543652 279016 543658
rect 278964 543594 279016 543600
rect 279068 543182 279096 660214
rect 279148 660204 279200 660210
rect 279148 660146 279200 660152
rect 279160 543250 279188 660146
rect 279240 660068 279292 660074
rect 279240 660010 279292 660016
rect 279252 543590 279280 660010
rect 279240 543584 279292 543590
rect 279240 543526 279292 543532
rect 279344 543318 279372 661710
rect 279436 543386 279464 663070
rect 279976 663060 280028 663066
rect 279976 663002 280028 663008
rect 279516 661564 279568 661570
rect 279516 661506 279568 661512
rect 279528 545902 279556 661506
rect 279608 660408 279660 660414
rect 279608 660350 279660 660356
rect 279516 545896 279568 545902
rect 279516 545838 279568 545844
rect 279620 545766 279648 660350
rect 279608 545760 279660 545766
rect 279608 545702 279660 545708
rect 279988 543522 280016 663002
rect 280068 661632 280120 661638
rect 280068 661574 280120 661580
rect 279976 543516 280028 543522
rect 279976 543458 280028 543464
rect 280080 543454 280108 661574
rect 296904 660000 296956 660006
rect 296904 659942 296956 659948
rect 296916 659841 296944 659942
rect 296902 659832 296958 659841
rect 296902 659767 296958 659776
rect 316144 654134 316172 683130
rect 317432 654134 317460 700334
rect 316144 654106 316724 654134
rect 317432 654106 317828 654134
rect 310428 642456 310480 642462
rect 310428 642398 310480 642404
rect 287612 642388 287664 642394
rect 287612 642330 287664 642336
rect 286508 642116 286560 642122
rect 286508 642058 286560 642064
rect 284208 641980 284260 641986
rect 284208 641922 284260 641928
rect 282734 641880 282790 641889
rect 282734 641815 282790 641824
rect 282748 639826 282776 641815
rect 284220 639962 284248 641922
rect 286520 639962 286548 642058
rect 287624 639962 287652 642330
rect 293132 642320 293184 642326
rect 293132 642262 293184 642268
rect 290924 641912 290976 641918
rect 290924 641854 290976 641860
rect 290936 639962 290964 641854
rect 293144 639962 293172 642262
rect 295248 642252 295300 642258
rect 295248 642194 295300 642200
rect 295260 639962 295288 642194
rect 300768 642184 300820 642190
rect 300768 642126 300820 642132
rect 296352 642048 296404 642054
rect 296352 641990 296404 641996
rect 296364 639962 296392 641990
rect 297548 641844 297600 641850
rect 297548 641786 297600 641792
rect 297560 639962 297588 641786
rect 300780 639962 300808 642126
rect 304170 641744 304226 641753
rect 304170 641679 304226 641688
rect 303068 640552 303120 640558
rect 303068 640494 303120 640500
rect 301962 640384 302018 640393
rect 301962 640319 302018 640328
rect 301976 639962 302004 640319
rect 303080 639962 303108 640494
rect 304184 639962 304212 641679
rect 310440 641034 310468 642398
rect 315856 641096 315908 641102
rect 315856 641038 315908 641044
rect 310428 641028 310480 641034
rect 310428 640970 310480 640976
rect 314108 641028 314160 641034
rect 314108 640970 314160 640976
rect 313004 640688 313056 640694
rect 313004 640630 313056 640636
rect 308588 640620 308640 640626
rect 308588 640562 308640 640568
rect 306194 640520 306250 640529
rect 306194 640455 306250 640464
rect 306208 639962 306236 640455
rect 308600 639962 308628 640562
rect 310336 640416 310388 640422
rect 310336 640358 310388 640364
rect 284004 639934 284248 639962
rect 286212 639934 286548 639962
rect 287316 639934 287652 639962
rect 290628 639934 290964 639962
rect 292836 639934 293172 639962
rect 295044 639934 295288 639962
rect 296148 639934 296392 639962
rect 297252 639934 297588 639962
rect 300564 639934 300808 639962
rect 301668 639934 302004 639962
rect 302772 639934 303108 639962
rect 303876 639934 304212 639962
rect 306084 639934 306236 639962
rect 308292 639934 308628 639962
rect 310348 639826 310376 640358
rect 311808 640348 311860 640354
rect 311808 640290 311860 640296
rect 311820 639962 311848 640290
rect 313016 639962 313044 640630
rect 314120 639962 314148 640970
rect 315212 640484 315264 640490
rect 315212 640426 315264 640432
rect 315224 639962 315252 640426
rect 311604 639934 311848 639962
rect 312708 639934 313044 639962
rect 313812 639934 314148 639962
rect 314916 639934 315252 639962
rect 315868 639826 315896 641038
rect 316696 639962 316724 654106
rect 317800 639962 317828 654106
rect 319444 641912 319496 641918
rect 319444 641854 319496 641860
rect 316696 639934 317124 639962
rect 317800 639934 318228 639962
rect 282748 639798 282900 639826
rect 310348 639798 310500 639826
rect 315868 639798 316020 639826
rect 299110 639432 299166 639441
rect 299166 639390 299460 639418
rect 319180 639402 319332 639418
rect 319168 639396 319332 639402
rect 299110 639367 299166 639376
rect 319220 639390 319332 639396
rect 319168 639338 319220 639344
rect 292028 639328 292080 639334
rect 282090 639296 282146 639305
rect 280172 639254 280692 639282
rect 281796 639254 282090 639282
rect 280172 551313 280200 639254
rect 285402 639296 285458 639305
rect 285108 639254 285402 639282
rect 282090 639231 282146 639240
rect 285402 639231 285458 639240
rect 288254 639296 288310 639305
rect 289634 639296 289690 639305
rect 288310 639254 288420 639282
rect 289524 639254 289634 639282
rect 288254 639231 288310 639240
rect 291732 639276 292028 639282
rect 294052 639328 294104 639334
rect 291732 639270 292080 639276
rect 293940 639276 294052 639282
rect 305092 639328 305144 639334
rect 298466 639296 298522 639305
rect 293940 639270 294104 639276
rect 291732 639254 292068 639270
rect 293940 639254 294092 639270
rect 298356 639254 298466 639282
rect 289634 639231 289690 639240
rect 304980 639276 305092 639282
rect 307484 639328 307536 639334
rect 304980 639270 305144 639276
rect 307188 639276 307484 639282
rect 309692 639328 309744 639334
rect 307188 639270 307536 639276
rect 309396 639276 309692 639282
rect 309396 639270 309744 639276
rect 304980 639254 305132 639270
rect 307188 639254 307524 639270
rect 309396 639254 309732 639270
rect 298466 639231 298522 639240
rect 301962 600672 302018 600681
rect 301668 600630 301962 600658
rect 303434 600672 303490 600681
rect 301962 600607 302018 600616
rect 302988 600630 303434 600658
rect 281552 600086 282348 600114
rect 282472 600086 282900 600114
rect 283024 600086 283452 600114
rect 283668 600086 284004 600114
rect 280158 551304 280214 551313
rect 280158 551239 280214 551248
rect 281552 547874 281580 600086
rect 282472 586514 282500 600086
rect 283024 599350 283052 600086
rect 283012 599344 283064 599350
rect 283012 599286 283064 599292
rect 282920 598188 282972 598194
rect 282920 598130 282972 598136
rect 281644 586486 282500 586514
rect 281644 573345 281672 586486
rect 281630 573336 281686 573345
rect 281630 573271 281686 573280
rect 282932 560969 282960 598130
rect 283024 570722 283052 599286
rect 283668 598194 283696 600086
rect 284542 599842 284570 600100
rect 284680 600086 285108 600114
rect 284542 599814 284616 599842
rect 284588 598262 284616 599814
rect 284576 598256 284628 598262
rect 284576 598198 284628 598204
rect 283656 598188 283708 598194
rect 283656 598130 283708 598136
rect 284680 586514 284708 600086
rect 285646 599842 285674 600100
rect 285600 599814 285674 599842
rect 285784 600086 286212 600114
rect 286764 600086 286916 600114
rect 285600 598194 285628 599814
rect 285588 598188 285640 598194
rect 285588 598130 285640 598136
rect 285784 586514 285812 600086
rect 286324 598188 286376 598194
rect 286324 598130 286376 598136
rect 284312 586486 284708 586514
rect 285692 586486 285812 586514
rect 284312 571985 284340 586486
rect 285692 583030 285720 586486
rect 285680 583024 285732 583030
rect 285680 582966 285732 582972
rect 286336 576162 286364 598130
rect 286888 597650 286916 600086
rect 287072 600086 287316 600114
rect 287440 600086 287868 600114
rect 288084 600086 288420 600114
rect 286876 597644 286928 597650
rect 286876 597586 286928 597592
rect 286324 576156 286376 576162
rect 286324 576098 286376 576104
rect 287072 574705 287100 600086
rect 287440 598210 287468 600086
rect 287164 598182 287468 598210
rect 287164 584458 287192 598182
rect 288084 594250 288112 600086
rect 288958 599842 288986 600100
rect 289096 600086 289524 600114
rect 290076 600086 290412 600114
rect 290628 600086 290964 600114
rect 288958 599814 289032 599842
rect 289004 598330 289032 599814
rect 288992 598324 289044 598330
rect 288992 598266 289044 598272
rect 289096 598210 289124 600086
rect 288452 598182 289124 598210
rect 288072 594244 288124 594250
rect 288072 594186 288124 594192
rect 288452 588606 288480 598182
rect 290384 597854 290412 600086
rect 290936 598398 290964 600086
rect 291166 599842 291194 600100
rect 291120 599814 291194 599842
rect 291304 600086 291732 600114
rect 291948 600086 292284 600114
rect 292684 600086 292836 600114
rect 292960 600086 293388 600114
rect 293604 600086 293940 600114
rect 290924 598392 290976 598398
rect 290924 598334 290976 598340
rect 291120 598194 291148 599814
rect 291108 598188 291160 598194
rect 291108 598130 291160 598136
rect 291200 598120 291252 598126
rect 291200 598062 291252 598068
rect 290372 597848 290424 597854
rect 290372 597790 290424 597796
rect 289084 597644 289136 597650
rect 289084 597586 289136 597592
rect 288440 588600 288492 588606
rect 288440 588542 288492 588548
rect 287152 584452 287204 584458
rect 287152 584394 287204 584400
rect 287058 574696 287114 574705
rect 287058 574631 287114 574640
rect 284298 571976 284354 571985
rect 284298 571911 284354 571920
rect 283012 570716 283064 570722
rect 283012 570658 283064 570664
rect 289096 560998 289124 597586
rect 289084 560992 289136 560998
rect 282918 560960 282974 560969
rect 289084 560934 289136 560940
rect 282918 560895 282974 560904
rect 291212 551342 291240 598062
rect 291304 595474 291332 600086
rect 291844 598188 291896 598194
rect 291844 598130 291896 598136
rect 291292 595468 291344 595474
rect 291292 595410 291344 595416
rect 291856 562358 291884 598130
rect 291948 598126 291976 600086
rect 292580 598188 292632 598194
rect 292580 598130 292632 598136
rect 291936 598120 291988 598126
rect 291936 598062 291988 598068
rect 292592 573374 292620 598130
rect 292684 574841 292712 600086
rect 292960 589966 292988 600086
rect 293604 598194 293632 600086
rect 294478 599842 294506 600100
rect 294616 600086 295044 600114
rect 295444 600086 295596 600114
rect 295812 600086 296148 600114
rect 296364 600086 296700 600114
rect 297252 600086 297588 600114
rect 297804 600086 298048 600114
rect 298356 600086 298692 600114
rect 298908 600086 299244 600114
rect 294478 599814 294552 599842
rect 294524 598534 294552 599814
rect 294512 598528 294564 598534
rect 294512 598470 294564 598476
rect 294616 598210 294644 600086
rect 293592 598188 293644 598194
rect 293592 598130 293644 598136
rect 293972 598182 294644 598210
rect 295340 598188 295392 598194
rect 293972 591326 294000 598182
rect 295340 598130 295392 598136
rect 294604 597848 294656 597854
rect 294604 597790 294656 597796
rect 293960 591320 294012 591326
rect 293960 591262 294012 591268
rect 292948 589960 293000 589966
rect 292948 589902 293000 589908
rect 292670 574832 292726 574841
rect 292670 574767 292726 574776
rect 292580 573368 292632 573374
rect 292580 573310 292632 573316
rect 294616 568041 294644 597790
rect 294602 568032 294658 568041
rect 294602 567967 294658 567976
rect 291844 562352 291896 562358
rect 291844 562294 291896 562300
rect 295352 551478 295380 598130
rect 295340 551472 295392 551478
rect 295340 551414 295392 551420
rect 295444 551410 295472 600086
rect 295812 598194 295840 600086
rect 295800 598188 295852 598194
rect 295800 598130 295852 598136
rect 296364 586514 296392 600086
rect 296720 599140 296772 599146
rect 296720 599082 296772 599088
rect 295536 586486 296392 586514
rect 295536 554062 295564 586486
rect 296732 565214 296760 599082
rect 297560 596834 297588 600086
rect 298020 599146 298048 600086
rect 298008 599140 298060 599146
rect 298008 599082 298060 599088
rect 298664 598806 298692 600086
rect 298652 598800 298704 598806
rect 298652 598742 298704 598748
rect 299216 598194 299244 600086
rect 299446 599842 299474 600100
rect 300012 600086 300348 600114
rect 300564 600086 300808 600114
rect 301116 600086 301452 600114
rect 299400 599814 299474 599842
rect 299400 598942 299428 599814
rect 300320 599010 300348 600086
rect 299480 599004 299532 599010
rect 299480 598946 299532 598952
rect 300308 599004 300360 599010
rect 300308 598946 300360 598952
rect 299388 598936 299440 598942
rect 299388 598878 299440 598884
rect 299388 598800 299440 598806
rect 299388 598742 299440 598748
rect 299204 598188 299256 598194
rect 299204 598130 299256 598136
rect 297548 596828 297600 596834
rect 297548 596770 297600 596776
rect 299400 580281 299428 598742
rect 299492 583001 299520 598946
rect 300124 598528 300176 598534
rect 300124 598470 300176 598476
rect 299478 582992 299534 583001
rect 299478 582927 299534 582936
rect 299386 580272 299442 580281
rect 299386 580207 299442 580216
rect 296720 565208 296772 565214
rect 296720 565150 296772 565156
rect 300136 563786 300164 598470
rect 300674 598224 300730 598233
rect 300674 598159 300676 598168
rect 300728 598159 300730 598168
rect 300676 598130 300728 598136
rect 300688 581641 300716 598130
rect 300780 598058 300808 600086
rect 300952 599888 301004 599894
rect 300952 599830 301004 599836
rect 300860 599412 300912 599418
rect 300860 599354 300912 599360
rect 300768 598052 300820 598058
rect 300768 597994 300820 598000
rect 300674 581632 300730 581641
rect 300674 581567 300730 581576
rect 300124 563780 300176 563786
rect 300124 563722 300176 563728
rect 300780 562426 300808 597994
rect 300872 577522 300900 599354
rect 300964 592657 300992 599830
rect 301424 599418 301452 600086
rect 302206 599894 302234 600100
rect 302772 600086 302924 600114
rect 302194 599888 302246 599894
rect 302194 599830 302246 599836
rect 302206 599706 302234 599830
rect 302160 599678 302234 599706
rect 301412 599412 301464 599418
rect 301412 599354 301464 599360
rect 302160 599214 302188 599678
rect 302148 599208 302200 599214
rect 302148 599150 302200 599156
rect 302238 598904 302294 598913
rect 302238 598839 302294 598848
rect 302252 595610 302280 598839
rect 302896 598194 302924 600086
rect 302988 598913 303016 600630
rect 306838 600672 306894 600681
rect 306636 600630 306838 600658
rect 303434 600607 303490 600616
rect 306838 600607 306894 600616
rect 307574 600672 307630 600681
rect 307574 600607 307630 600616
rect 305932 600222 306084 600250
rect 303876 600086 304212 600114
rect 304428 600086 304764 600114
rect 302974 598904 303030 598913
rect 302974 598839 303030 598848
rect 304184 598670 304212 600086
rect 304736 598874 304764 600086
rect 304966 599842 304994 600100
rect 305532 600086 305868 600114
rect 304920 599814 304994 599842
rect 304724 598868 304776 598874
rect 304724 598810 304776 598816
rect 304172 598664 304224 598670
rect 304172 598606 304224 598612
rect 304632 598664 304684 598670
rect 304632 598606 304684 598612
rect 302884 598188 302936 598194
rect 302884 598130 302936 598136
rect 304644 596174 304672 598606
rect 304736 598346 304764 598810
rect 304920 598602 304948 599814
rect 305000 599276 305052 599282
rect 305000 599218 305052 599224
rect 304908 598596 304960 598602
rect 304908 598538 304960 598544
rect 304736 598318 304856 598346
rect 304644 596146 304764 596174
rect 302240 595604 302292 595610
rect 302240 595546 302292 595552
rect 300950 592648 301006 592657
rect 300950 592583 301006 592592
rect 300860 577516 300912 577522
rect 300860 577458 300912 577464
rect 304736 570654 304764 596146
rect 304724 570648 304776 570654
rect 304724 570590 304776 570596
rect 300768 562420 300820 562426
rect 300768 562362 300820 562368
rect 304828 561066 304856 598318
rect 304816 561060 304868 561066
rect 304816 561002 304868 561008
rect 295524 554056 295576 554062
rect 295524 553998 295576 554004
rect 295432 551404 295484 551410
rect 295432 551346 295484 551352
rect 291200 551336 291252 551342
rect 291200 551278 291252 551284
rect 304920 548554 304948 598538
rect 305012 566506 305040 599218
rect 305840 598738 305868 600086
rect 305932 599282 305960 600222
rect 306760 600086 307188 600114
rect 306380 599888 306432 599894
rect 306380 599830 306432 599836
rect 305920 599276 305972 599282
rect 305920 599218 305972 599224
rect 305828 598732 305880 598738
rect 305828 598674 305880 598680
rect 306288 598732 306340 598738
rect 306288 598674 306340 598680
rect 305000 566500 305052 566506
rect 305000 566442 305052 566448
rect 304908 548548 304960 548554
rect 304908 548490 304960 548496
rect 281540 547868 281592 547874
rect 281540 547810 281592 547816
rect 297456 543652 297508 543658
rect 297456 543594 297508 543600
rect 280068 543448 280120 543454
rect 280068 543390 280120 543396
rect 296166 543416 296222 543425
rect 279424 543380 279476 543386
rect 296166 543351 296222 543360
rect 279424 543322 279476 543328
rect 279332 543312 279384 543318
rect 279332 543254 279384 543260
rect 279148 543244 279200 543250
rect 279148 543186 279200 543192
rect 279056 543176 279108 543182
rect 279056 543118 279108 543124
rect 278136 543108 278188 543114
rect 278136 543050 278188 543056
rect 296180 542745 296208 543351
rect 279790 542736 279846 542745
rect 279790 542671 279846 542680
rect 292578 542736 292634 542745
rect 292578 542671 292634 542680
rect 296166 542736 296222 542745
rect 296166 542671 296222 542680
rect 279700 542632 279752 542638
rect 279700 542574 279752 542580
rect 279608 542564 279660 542570
rect 279608 542506 279660 542512
rect 279516 542428 279568 542434
rect 279516 542370 279568 542376
rect 278320 539708 278372 539714
rect 278320 539650 278372 539656
rect 278136 534132 278188 534138
rect 278136 534074 278188 534080
rect 278044 137964 278096 137970
rect 278044 137906 278096 137912
rect 278148 64870 278176 534074
rect 278228 447160 278280 447166
rect 278228 447102 278280 447108
rect 278240 114510 278268 447102
rect 278332 281110 278360 539650
rect 278780 496188 278832 496194
rect 278780 496130 278832 496136
rect 278320 281104 278372 281110
rect 278320 281046 278372 281052
rect 278228 114504 278280 114510
rect 278228 114446 278280 114452
rect 278136 64864 278188 64870
rect 278136 64806 278188 64812
rect 278792 16574 278820 496130
rect 279424 488572 279476 488578
rect 279424 488514 279476 488520
rect 279436 125594 279464 488514
rect 279528 279954 279556 542370
rect 279516 279948 279568 279954
rect 279516 279890 279568 279896
rect 279620 279886 279648 542506
rect 279712 280022 279740 542574
rect 279804 281314 279832 542671
rect 279884 542496 279936 542502
rect 279884 542438 279936 542444
rect 279896 281926 279924 542438
rect 292592 540138 292620 542671
rect 294512 542632 294564 542638
rect 294512 542574 294564 542580
rect 293960 542564 294012 542570
rect 293960 542506 294012 542512
rect 292592 540110 292666 540138
rect 292638 539852 292666 540110
rect 293972 539866 294000 542506
rect 294524 539866 294552 542574
rect 295340 542496 295392 542502
rect 295340 542438 295392 542444
rect 297178 542464 297234 542473
rect 295352 539866 295380 542438
rect 295984 542428 296036 542434
rect 297178 542399 297234 542408
rect 295984 542370 296036 542376
rect 295996 539866 296024 542370
rect 293972 539838 294124 539866
rect 294524 539838 294860 539866
rect 295352 539838 295596 539866
rect 295996 539838 296332 539866
rect 287886 539744 287942 539753
rect 283484 539714 283820 539730
rect 283472 539708 283820 539714
rect 283524 539702 283820 539708
rect 297192 539730 297220 542399
rect 297468 539866 297496 543594
rect 300400 543584 300452 543590
rect 300400 543526 300452 543532
rect 298190 542872 298246 542881
rect 298190 542807 298246 542816
rect 298204 539866 298232 542807
rect 298926 542600 298982 542609
rect 298926 542535 298982 542544
rect 298940 539866 298968 542535
rect 299938 542464 299994 542473
rect 299938 542399 299994 542408
rect 299952 540138 299980 542399
rect 299952 540110 300026 540138
rect 297468 539838 297804 539866
rect 298204 539838 298540 539866
rect 298940 539838 299276 539866
rect 299998 539852 300026 540110
rect 300412 539866 300440 543526
rect 301136 543516 301188 543522
rect 301136 543458 301188 543464
rect 301148 539866 301176 543458
rect 302608 543448 302660 543454
rect 302608 543390 302660 543396
rect 301870 543144 301926 543153
rect 301870 543079 301926 543088
rect 301884 539866 301912 543079
rect 302620 539866 302648 543390
rect 303804 543380 303856 543386
rect 303804 543322 303856 543328
rect 300412 539838 300748 539866
rect 301148 539838 301484 539866
rect 301884 539838 302220 539866
rect 302620 539838 302956 539866
rect 287942 539702 288236 539730
rect 297068 539702 297220 539730
rect 287886 539679 287942 539688
rect 283472 539650 283524 539656
rect 286416 539640 286468 539646
rect 283378 539608 283434 539617
rect 280804 539572 280856 539578
rect 280804 539514 280856 539520
rect 281000 539566 282348 539594
rect 283084 539566 283378 539594
rect 279884 281920 279936 281926
rect 279884 281862 279936 281868
rect 279792 281308 279844 281314
rect 279792 281250 279844 281256
rect 280816 281178 280844 539514
rect 281000 281246 281028 539566
rect 286138 539608 286194 539617
rect 284220 539578 284556 539594
rect 283378 539543 283434 539552
rect 284208 539572 284556 539578
rect 284260 539566 284556 539572
rect 284956 539566 285292 539594
rect 286028 539566 286138 539594
rect 284208 539514 284260 539520
rect 284956 539510 284984 539566
rect 287610 539608 287666 539617
rect 286468 539588 286764 539594
rect 286416 539582 286764 539588
rect 286428 539566 286764 539582
rect 287500 539566 287610 539594
rect 286138 539543 286194 539552
rect 287610 539543 287666 539552
rect 288622 539608 288678 539617
rect 289358 539608 289414 539617
rect 288678 539566 288972 539594
rect 288622 539543 288678 539552
rect 290554 539608 290610 539617
rect 289414 539566 289708 539594
rect 290444 539566 290554 539594
rect 289358 539543 289414 539552
rect 290554 539543 290610 539552
rect 290830 539608 290886 539617
rect 291566 539608 291622 539617
rect 290886 539566 291180 539594
rect 290830 539543 290886 539552
rect 293038 539608 293094 539617
rect 291622 539566 291916 539594
rect 291566 539543 291622 539552
rect 303816 539594 303844 543322
rect 305552 543312 305604 543318
rect 305552 543254 305604 543260
rect 304078 542872 304134 542881
rect 304078 542807 304134 542816
rect 304092 539866 304120 542807
rect 304998 542736 305054 542745
rect 304998 542671 305054 542680
rect 305012 539866 305040 542671
rect 305564 539866 305592 543254
rect 306300 541754 306328 598674
rect 306392 572014 306420 599830
rect 306760 590034 306788 600086
rect 307588 596174 307616 600607
rect 307726 599894 307754 600100
rect 307714 599888 307766 599894
rect 307714 599830 307766 599836
rect 308278 599842 308306 600100
rect 308416 600086 308844 600114
rect 309244 600086 309396 600114
rect 309520 600086 309948 600114
rect 310164 600086 310500 600114
rect 310624 600086 311052 600114
rect 311176 600086 311604 600114
rect 308278 599814 308352 599842
rect 308324 598534 308352 599814
rect 308312 598528 308364 598534
rect 308312 598470 308364 598476
rect 307588 596146 307708 596174
rect 306748 590028 306800 590034
rect 306748 589970 306800 589976
rect 306380 572008 306432 572014
rect 306380 571950 306432 571956
rect 307680 545086 307708 596146
rect 308416 586514 308444 600086
rect 309140 598120 309192 598126
rect 309140 598062 309192 598068
rect 307772 586486 308444 586514
rect 307772 584526 307800 586486
rect 307760 584520 307812 584526
rect 307760 584462 307812 584468
rect 307668 545080 307720 545086
rect 307668 545022 307720 545028
rect 307022 543280 307078 543289
rect 307022 543215 307078 543224
rect 306378 542464 306434 542473
rect 306378 542399 306434 542408
rect 306288 541748 306340 541754
rect 306288 541690 306340 541696
rect 306392 539866 306420 542399
rect 307036 539866 307064 543215
rect 308494 542600 308550 542609
rect 308494 542535 308550 542544
rect 308402 542464 308458 542473
rect 308402 542399 308458 542408
rect 308416 539866 308444 542399
rect 304092 539838 304428 539866
rect 305012 539838 305164 539866
rect 305564 539838 305900 539866
rect 306392 539838 306636 539866
rect 307036 539838 307372 539866
rect 308108 539838 308444 539866
rect 308508 539866 308536 542535
rect 309152 541686 309180 598062
rect 309244 552838 309272 600086
rect 309520 586514 309548 600086
rect 310164 598126 310192 600086
rect 310152 598120 310204 598126
rect 310624 598108 310652 600086
rect 311072 598188 311124 598194
rect 311072 598130 311124 598136
rect 310152 598062 310204 598068
rect 310532 598080 310652 598108
rect 309336 586486 309548 586514
rect 309336 563825 309364 586486
rect 310532 580310 310560 598080
rect 311084 596902 311112 598130
rect 311072 596896 311124 596902
rect 311072 596838 311124 596844
rect 311176 594114 311204 600086
rect 312142 599842 312170 600100
rect 312096 599814 312170 599842
rect 312372 600086 312708 600114
rect 312924 600086 313260 600114
rect 313384 600086 313812 600114
rect 314028 600086 314364 600114
rect 314764 600086 314916 600114
rect 315132 600086 315468 600114
rect 315684 600086 316020 600114
rect 316572 600086 316908 600114
rect 317124 600086 317368 600114
rect 311992 598188 312044 598194
rect 311992 598130 312044 598136
rect 311900 598120 311952 598126
rect 311900 598062 311952 598068
rect 311164 594108 311216 594114
rect 311164 594050 311216 594056
rect 310520 580304 310572 580310
rect 310520 580246 310572 580252
rect 311912 568177 311940 598062
rect 312004 588674 312032 598130
rect 312096 592006 312124 599814
rect 312372 598126 312400 600086
rect 312924 598194 312952 600086
rect 312912 598188 312964 598194
rect 312912 598130 312964 598136
rect 313280 598188 313332 598194
rect 313280 598130 313332 598136
rect 312360 598120 312412 598126
rect 312360 598062 312412 598068
rect 312084 592000 312136 592006
rect 312084 591942 312136 591948
rect 311992 588668 312044 588674
rect 311992 588610 312044 588616
rect 311898 568168 311954 568177
rect 311898 568103 311954 568112
rect 309322 563816 309378 563825
rect 309322 563751 309378 563760
rect 309232 552832 309284 552838
rect 309232 552774 309284 552780
rect 313292 545766 313320 598130
rect 313384 573442 313412 600086
rect 314028 598194 314056 600086
rect 314016 598188 314068 598194
rect 314016 598130 314068 598136
rect 314660 598188 314712 598194
rect 314660 598130 314712 598136
rect 313372 573436 313424 573442
rect 313372 573378 313424 573384
rect 314672 558249 314700 598130
rect 314764 569294 314792 600086
rect 315132 598194 315160 600086
rect 315120 598188 315172 598194
rect 315120 598130 315172 598136
rect 315684 586514 315712 600086
rect 316880 598194 316908 600086
rect 317340 598466 317368 600086
rect 317432 600086 317676 600114
rect 317328 598460 317380 598466
rect 317328 598402 317380 598408
rect 316868 598188 316920 598194
rect 316868 598130 316920 598136
rect 316684 592000 316736 592006
rect 316684 591942 316736 591948
rect 314856 586486 315712 586514
rect 314856 576230 314884 586486
rect 314844 576224 314896 576230
rect 314844 576166 314896 576172
rect 314752 569288 314804 569294
rect 314752 569230 314804 569236
rect 314658 558240 314714 558249
rect 314658 558175 314714 558184
rect 316696 546446 316724 591942
rect 316684 546440 316736 546446
rect 316684 546382 316736 546388
rect 313648 545896 313700 545902
rect 313648 545838 313700 545844
rect 312912 545760 312964 545766
rect 312912 545702 312964 545708
rect 313280 545760 313332 545766
rect 313280 545702 313332 545708
rect 312266 542872 312322 542881
rect 312266 542807 312322 542816
rect 310702 542736 310758 542745
rect 310702 542671 310758 542680
rect 309966 542600 310022 542609
rect 309966 542535 310022 542544
rect 309414 542464 309470 542473
rect 309414 542399 309470 542408
rect 309140 541680 309192 541686
rect 309140 541622 309192 541628
rect 309428 539866 309456 542399
rect 309980 539866 310008 542535
rect 310716 539866 310744 542671
rect 311438 542464 311494 542473
rect 311438 542399 311494 542408
rect 311452 539866 311480 542399
rect 312280 539866 312308 542807
rect 312924 539866 312952 545702
rect 313660 539866 313688 545838
rect 316040 543244 316092 543250
rect 316040 543186 316092 543192
rect 315120 543176 315172 543182
rect 315120 543118 315172 543124
rect 314844 543040 314896 543046
rect 314844 542982 314896 542988
rect 308508 539838 308844 539866
rect 309428 539838 309580 539866
rect 309980 539838 310316 539866
rect 310716 539838 311052 539866
rect 311452 539838 311788 539866
rect 312280 539838 312524 539866
rect 312924 539838 313260 539866
rect 313660 539838 313996 539866
rect 314856 539594 314884 542982
rect 315132 539866 315160 543118
rect 315132 539838 315468 539866
rect 316052 539730 316080 543186
rect 316592 543108 316644 543114
rect 316592 543050 316644 543056
rect 316604 539866 316632 543050
rect 317432 540258 317460 600086
rect 319456 566409 319484 641854
rect 320824 640416 320876 640422
rect 320824 640358 320876 640364
rect 319720 639532 319772 639538
rect 319720 639474 319772 639480
rect 319536 639464 319588 639470
rect 319536 639406 319588 639412
rect 319548 598058 319576 639406
rect 319732 625154 319760 639474
rect 319640 625126 319760 625154
rect 319640 598233 319668 625126
rect 319626 598224 319682 598233
rect 319626 598159 319682 598168
rect 319536 598052 319588 598058
rect 319536 597994 319588 598000
rect 319442 566400 319498 566409
rect 319442 566335 319498 566344
rect 320180 563712 320232 563718
rect 320180 563654 320232 563660
rect 317510 543688 317566 543697
rect 317510 543623 317566 543632
rect 317420 540252 317472 540258
rect 317420 540194 317472 540200
rect 316604 539838 316940 539866
rect 316052 539702 316204 539730
rect 293094 539566 293388 539594
rect 303692 539566 303844 539594
rect 314732 539566 314884 539594
rect 317524 539594 317552 543623
rect 317524 539566 317676 539594
rect 293038 539543 293094 539552
rect 281172 539504 281224 539510
rect 281172 539446 281224 539452
rect 284944 539504 284996 539510
rect 284944 539446 284996 539452
rect 281184 281382 281212 539446
rect 320192 537538 320220 563654
rect 320180 537532 320232 537538
rect 320180 537474 320232 537480
rect 320192 537373 320220 537474
rect 320178 537364 320234 537373
rect 320178 537299 320234 537308
rect 320364 513324 320416 513330
rect 320364 513266 320416 513272
rect 320376 512213 320404 513266
rect 320362 512204 320418 512213
rect 320362 512139 320418 512148
rect 320364 510876 320416 510882
rect 320362 510844 320364 510853
rect 320640 510876 320692 510882
rect 320416 510844 320418 510853
rect 320640 510818 320692 510824
rect 320362 510779 320418 510788
rect 320088 510604 320140 510610
rect 320088 510546 320140 510552
rect 320100 510173 320128 510546
rect 320456 510536 320508 510542
rect 320456 510478 320508 510484
rect 320086 510164 320142 510173
rect 320086 510099 320142 510108
rect 319350 509960 319406 509969
rect 319350 509895 319406 509904
rect 319364 509234 319392 509895
rect 320468 509561 320496 510478
rect 320454 509552 320510 509561
rect 320454 509487 320510 509496
rect 319180 509206 319392 509234
rect 320180 509244 320232 509250
rect 319076 508292 319128 508298
rect 319076 508234 319128 508240
rect 319088 507890 319116 508234
rect 319076 507884 319128 507890
rect 319076 507826 319128 507832
rect 318984 506524 319036 506530
rect 318984 506466 319036 506472
rect 318892 505572 318944 505578
rect 318892 505514 318944 505520
rect 296628 500404 296680 500410
rect 296628 500346 296680 500352
rect 295248 500336 295300 500342
rect 295248 500278 295300 500284
rect 292764 500268 292816 500274
rect 292764 500210 292816 500216
rect 281552 500126 282348 500154
rect 281552 324290 281580 500126
rect 283070 499882 283098 500140
rect 283208 500126 283820 500154
rect 283070 499854 283144 499882
rect 282184 498840 282236 498846
rect 282184 498782 282236 498788
rect 281540 324284 281592 324290
rect 281540 324226 281592 324232
rect 281172 281376 281224 281382
rect 281172 281318 281224 281324
rect 280988 281240 281040 281246
rect 280988 281182 281040 281188
rect 280804 281172 280856 281178
rect 280804 281114 280856 281120
rect 279700 280016 279752 280022
rect 279700 279958 279752 279964
rect 279608 279880 279660 279886
rect 279608 279822 279660 279828
rect 279424 125588 279476 125594
rect 279424 125530 279476 125536
rect 282196 67590 282224 498782
rect 282920 345704 282972 345710
rect 282920 345646 282972 345652
rect 282184 67584 282236 67590
rect 282184 67526 282236 67532
rect 282932 16574 282960 345646
rect 283116 342922 283144 499854
rect 283104 342916 283156 342922
rect 283104 342858 283156 342864
rect 283208 227118 283236 500126
rect 284542 499882 284570 500140
rect 284680 500126 285292 500154
rect 285876 500126 286028 500154
rect 286428 500126 286764 500154
rect 287164 500126 287500 500154
rect 287900 500126 288236 500154
rect 288544 500126 288972 500154
rect 289372 500126 289708 500154
rect 284542 499854 284616 499882
rect 284588 496874 284616 499854
rect 284576 496868 284628 496874
rect 284576 496810 284628 496816
rect 284680 489914 284708 500126
rect 285680 494760 285732 494766
rect 285680 494702 285732 494708
rect 284312 489886 284708 489914
rect 284312 330546 284340 489886
rect 284944 452668 284996 452674
rect 284944 452610 284996 452616
rect 284300 330540 284352 330546
rect 284300 330482 284352 330488
rect 283196 227112 283248 227118
rect 283196 227054 283248 227060
rect 284956 117298 284984 452610
rect 285128 332240 285180 332246
rect 285128 332182 285180 332188
rect 285036 329928 285088 329934
rect 285036 329870 285088 329876
rect 285048 317422 285076 329870
rect 285140 320142 285168 332182
rect 285128 320136 285180 320142
rect 285128 320078 285180 320084
rect 285036 317416 285088 317422
rect 285036 317358 285088 317364
rect 285036 295384 285088 295390
rect 285036 295326 285088 295332
rect 285048 281382 285076 295326
rect 285036 281376 285088 281382
rect 285036 281318 285088 281324
rect 284944 117292 284996 117298
rect 284944 117234 284996 117240
rect 285692 16574 285720 494702
rect 285876 491978 285904 500126
rect 286428 499574 286456 500126
rect 286244 499546 286456 499574
rect 285864 491972 285916 491978
rect 285864 491914 285916 491920
rect 286244 489914 286272 499546
rect 286324 496868 286376 496874
rect 286324 496810 286376 496816
rect 285784 489886 286272 489914
rect 285784 341562 285812 489886
rect 285772 341556 285824 341562
rect 285772 341498 285824 341504
rect 286336 333334 286364 496810
rect 287060 494692 287112 494698
rect 287060 494634 287112 494640
rect 286324 333328 286376 333334
rect 286324 333270 286376 333276
rect 286324 330540 286376 330546
rect 286324 330482 286376 330488
rect 286336 292534 286364 330482
rect 286324 292528 286376 292534
rect 286324 292470 286376 292476
rect 287072 278254 287100 494634
rect 287164 352578 287192 500126
rect 287900 494698 287928 500126
rect 287888 494692 287940 494698
rect 287888 494634 287940 494640
rect 288440 494692 288492 494698
rect 288440 494634 288492 494640
rect 287704 418192 287756 418198
rect 287704 418134 287756 418140
rect 287152 352572 287204 352578
rect 287152 352514 287204 352520
rect 287716 279002 287744 418134
rect 287796 365764 287848 365770
rect 287796 365706 287848 365712
rect 287808 318782 287836 365706
rect 288452 347070 288480 494634
rect 288544 354006 288572 500126
rect 289372 494698 289400 500126
rect 290430 499882 290458 500140
rect 290568 500126 291180 500154
rect 291304 500126 291916 500154
rect 290430 499854 290504 499882
rect 290476 497826 290504 499854
rect 290464 497820 290516 497826
rect 290464 497762 290516 497768
rect 289360 494692 289412 494698
rect 289360 494634 289412 494640
rect 290568 489914 290596 500126
rect 289924 489886 290596 489914
rect 289084 465112 289136 465118
rect 289084 465054 289136 465060
rect 288532 354000 288584 354006
rect 288532 353942 288584 353948
rect 288440 347064 288492 347070
rect 288440 347006 288492 347012
rect 287796 318776 287848 318782
rect 287796 318718 287848 318724
rect 287704 278996 287756 279002
rect 287704 278938 287756 278944
rect 287060 278248 287112 278254
rect 287060 278190 287112 278196
rect 287704 201544 287756 201550
rect 287704 201486 287756 201492
rect 287716 87650 287744 201486
rect 289096 120086 289124 465054
rect 289176 382288 289228 382294
rect 289176 382230 289228 382236
rect 289188 285666 289216 382230
rect 289268 353320 289320 353326
rect 289268 353262 289320 353268
rect 289176 285660 289228 285666
rect 289176 285602 289228 285608
rect 289280 279070 289308 353262
rect 289820 351212 289872 351218
rect 289820 351154 289872 351160
rect 289268 279064 289320 279070
rect 289268 279006 289320 279012
rect 289084 120080 289136 120086
rect 289084 120022 289136 120028
rect 287704 87644 287756 87650
rect 287704 87586 287756 87592
rect 278792 16546 279096 16574
rect 282932 16546 283144 16574
rect 285692 16546 286640 16574
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 283116 480 283144 16546
rect 286612 480 286640 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 354 289860 351154
rect 289924 338774 289952 489886
rect 289912 338768 289964 338774
rect 289912 338710 289964 338716
rect 291304 334626 291332 500126
rect 292638 499882 292666 500140
rect 292592 499854 292666 499882
rect 291936 497888 291988 497894
rect 291936 497830 291988 497836
rect 291844 434784 291896 434790
rect 291844 434726 291896 434732
rect 291292 334620 291344 334626
rect 291292 334562 291344 334568
rect 291856 88330 291884 434726
rect 291948 220250 291976 497830
rect 292028 491972 292080 491978
rect 292028 491914 292080 491920
rect 292040 288386 292068 491914
rect 292120 331560 292172 331566
rect 292120 331502 292172 331508
rect 292132 325650 292160 331502
rect 292120 325644 292172 325650
rect 292120 325586 292172 325592
rect 292592 303210 292620 499854
rect 292580 303204 292632 303210
rect 292580 303146 292632 303152
rect 292028 288380 292080 288386
rect 292028 288322 292080 288328
rect 291936 220244 291988 220250
rect 291936 220186 291988 220192
rect 291844 88324 291896 88330
rect 291844 88266 291896 88272
rect 292776 16574 292804 500210
rect 292868 500126 293388 500154
rect 292868 313274 292896 500126
rect 294110 499882 294138 500140
rect 294248 500126 294860 500154
rect 294110 499854 294184 499882
rect 294156 496738 294184 499854
rect 294144 496732 294196 496738
rect 294144 496674 294196 496680
rect 294248 489914 294276 500126
rect 294604 497956 294656 497962
rect 294604 497898 294656 497904
rect 293972 489886 294276 489914
rect 293222 332208 293278 332217
rect 293222 332143 293278 332152
rect 292856 313268 292908 313274
rect 292856 313210 292908 313216
rect 293236 218754 293264 332143
rect 293868 331764 293920 331770
rect 293868 331706 293920 331712
rect 293406 331528 293462 331537
rect 293406 331463 293462 331472
rect 293316 306400 293368 306406
rect 293316 306342 293368 306348
rect 293328 278798 293356 306342
rect 293316 278792 293368 278798
rect 293316 278734 293368 278740
rect 293420 227050 293448 331463
rect 293776 331424 293828 331430
rect 293776 331366 293828 331372
rect 293684 331288 293736 331294
rect 293684 331230 293736 331236
rect 293408 227044 293460 227050
rect 293408 226986 293460 226992
rect 293696 222902 293724 331230
rect 293788 222970 293816 331366
rect 293880 223038 293908 331706
rect 293972 303550 294000 489886
rect 293960 303544 294012 303550
rect 293960 303486 294012 303492
rect 293868 223032 293920 223038
rect 293868 222974 293920 222980
rect 293776 222964 293828 222970
rect 293776 222906 293828 222912
rect 293684 222896 293736 222902
rect 293684 222838 293736 222844
rect 294616 220182 294644 497898
rect 295156 332104 295208 332110
rect 295156 332046 295208 332052
rect 294972 331968 295024 331974
rect 294972 331910 295024 331916
rect 294696 303204 294748 303210
rect 294696 303146 294748 303152
rect 294708 278390 294736 303146
rect 294788 300892 294840 300898
rect 294788 300834 294840 300840
rect 294800 278866 294828 300834
rect 294788 278860 294840 278866
rect 294788 278802 294840 278808
rect 294984 278458 295012 331910
rect 295064 331900 295116 331906
rect 295064 331842 295116 331848
rect 295076 278730 295104 331842
rect 295064 278724 295116 278730
rect 295064 278666 295116 278672
rect 294972 278452 295024 278458
rect 294972 278394 295024 278400
rect 294696 278384 294748 278390
rect 294696 278326 294748 278332
rect 295168 278322 295196 332046
rect 295156 278316 295208 278322
rect 295156 278258 295208 278264
rect 294604 220176 294656 220182
rect 294604 220118 294656 220124
rect 293224 218748 293276 218754
rect 293224 218690 293276 218696
rect 295260 60178 295288 500278
rect 295352 500126 295596 500154
rect 295904 500126 296332 500154
rect 295352 278526 295380 500126
rect 295904 489914 295932 500126
rect 296074 498808 296130 498817
rect 296074 498743 296130 498752
rect 295984 496732 296036 496738
rect 295984 496674 296036 496680
rect 295444 489886 295932 489914
rect 295444 289678 295472 489886
rect 295432 289672 295484 289678
rect 295432 289614 295484 289620
rect 295430 282160 295486 282169
rect 295430 282095 295486 282104
rect 295444 282062 295472 282095
rect 295432 282056 295484 282062
rect 295432 281998 295484 282004
rect 295340 278520 295392 278526
rect 295340 278462 295392 278468
rect 295996 278186 296024 496674
rect 296088 281994 296116 498743
rect 296536 497480 296588 497486
rect 296536 497422 296588 497428
rect 296168 342304 296220 342310
rect 296168 342246 296220 342252
rect 296076 281988 296128 281994
rect 296076 281930 296128 281936
rect 296180 278934 296208 342246
rect 296444 332172 296496 332178
rect 296444 332114 296496 332120
rect 296352 332036 296404 332042
rect 296352 331978 296404 331984
rect 296260 331628 296312 331634
rect 296260 331570 296312 331576
rect 296272 279546 296300 331570
rect 296260 279540 296312 279546
rect 296260 279482 296312 279488
rect 296168 278928 296220 278934
rect 296168 278870 296220 278876
rect 296364 278662 296392 331978
rect 296352 278656 296404 278662
rect 296352 278598 296404 278604
rect 296456 278594 296484 332114
rect 296548 331945 296576 497422
rect 296534 331936 296590 331945
rect 296534 331871 296590 331880
rect 296534 331800 296590 331809
rect 296534 331735 296590 331744
rect 296444 278588 296496 278594
rect 296444 278530 296496 278536
rect 295984 278180 296036 278186
rect 295984 278122 296036 278128
rect 295982 204232 296038 204241
rect 295982 204167 296038 204176
rect 295996 91798 296024 204167
rect 295984 91792 296036 91798
rect 295984 91734 296036 91740
rect 295248 60172 295300 60178
rect 295248 60114 295300 60120
rect 292776 16546 293264 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 296548 3806 296576 331735
rect 296640 60246 296668 500346
rect 296824 500126 297068 500154
rect 297468 500126 297804 500154
rect 298112 500126 298540 500154
rect 298848 500126 299276 500154
rect 299676 500126 300012 500154
rect 300412 500126 300748 500154
rect 300964 500126 301484 500154
rect 301884 500126 302220 500154
rect 302436 500126 302956 500154
rect 296720 493468 296772 493474
rect 296720 493410 296772 493416
rect 296732 340202 296760 493410
rect 296824 341698 296852 500126
rect 297468 493474 297496 500126
rect 297456 493468 297508 493474
rect 297456 493410 297508 493416
rect 297640 460216 297692 460222
rect 297640 460158 297692 460164
rect 296812 341692 296864 341698
rect 296812 341634 296864 341640
rect 296720 340196 296772 340202
rect 296720 340138 296772 340144
rect 297362 329760 297418 329769
rect 297362 329695 297418 329704
rect 297270 325000 297326 325009
rect 297270 324935 297326 324944
rect 297086 320240 297142 320249
rect 297086 320175 297142 320184
rect 296994 301200 297050 301209
rect 296994 301135 297050 301144
rect 296810 217696 296866 217705
rect 296810 217631 296866 217640
rect 296824 216714 296852 217631
rect 296812 216708 296864 216714
rect 296812 216650 296864 216656
rect 296810 202736 296866 202745
rect 296810 202671 296866 202680
rect 296824 201550 296852 202671
rect 296812 201544 296864 201550
rect 296812 201486 296864 201492
rect 296810 166832 296866 166841
rect 296810 166767 296866 166776
rect 296824 165646 296852 166767
rect 296812 165640 296864 165646
rect 296812 165582 296864 165588
rect 296810 157856 296866 157865
rect 296810 157791 296866 157800
rect 296824 157418 296852 157791
rect 296812 157412 296864 157418
rect 296812 157354 296864 157360
rect 296810 148880 296866 148889
rect 296810 148815 296866 148824
rect 296824 147694 296852 148815
rect 296812 147688 296864 147694
rect 296812 147630 296864 147636
rect 296812 136604 296864 136610
rect 296812 136546 296864 136552
rect 296824 135425 296852 136546
rect 296810 135416 296866 135425
rect 296810 135351 296866 135360
rect 296812 118652 296864 118658
rect 296812 118594 296864 118600
rect 296824 117473 296852 118594
rect 296810 117464 296866 117473
rect 296810 117399 296866 117408
rect 297008 102513 297036 301135
rect 296994 102504 297050 102513
rect 296994 102439 297050 102448
rect 297100 92041 297128 320175
rect 297178 318880 297234 318889
rect 297178 318815 297234 318824
rect 297192 275398 297220 318815
rect 297284 316062 297312 324935
rect 297272 316056 297324 316062
rect 297272 315998 297324 316004
rect 297376 279478 297404 329695
rect 297454 328400 297510 328409
rect 297454 328335 297510 328344
rect 297364 279472 297416 279478
rect 297364 279414 297416 279420
rect 297468 276758 297496 328335
rect 297546 326360 297602 326369
rect 297546 326295 297602 326304
rect 297456 276752 297508 276758
rect 297456 276694 297508 276700
rect 297180 275392 297232 275398
rect 297180 275334 297232 275340
rect 297560 273970 297588 326295
rect 297652 284209 297680 460158
rect 297824 344412 297876 344418
rect 297824 344354 297876 344360
rect 297732 324284 297784 324290
rect 297732 324226 297784 324232
rect 297744 323649 297772 324226
rect 297730 323640 297786 323649
rect 297730 323575 297786 323584
rect 297732 318776 297784 318782
rect 297732 318718 297784 318724
rect 297744 317529 297772 318718
rect 297730 317520 297786 317529
rect 297730 317455 297786 317464
rect 297732 317416 297784 317422
rect 297732 317358 297784 317364
rect 297744 316169 297772 317358
rect 297730 316160 297786 316169
rect 297730 316095 297786 316104
rect 297732 316056 297784 316062
rect 297732 315998 297784 316004
rect 297744 296714 297772 315998
rect 297836 299169 297864 344354
rect 298112 333384 298140 500126
rect 298848 492658 298876 500126
rect 299480 494692 299532 494698
rect 299480 494634 299532 494640
rect 298836 492652 298888 492658
rect 298836 492594 298888 492600
rect 299020 348424 299072 348430
rect 299020 348366 299072 348372
rect 298560 334756 298612 334762
rect 298560 334698 298612 334704
rect 297928 333356 298140 333384
rect 297928 314809 297956 333356
rect 298008 333260 298060 333266
rect 298008 333202 298060 333208
rect 297914 314800 297970 314809
rect 297914 314735 297970 314744
rect 297916 313268 297968 313274
rect 297916 313210 297968 313216
rect 297928 312769 297956 313210
rect 297914 312760 297970 312769
rect 297914 312695 297970 312704
rect 298020 311409 298048 333202
rect 298006 311400 298062 311409
rect 298006 311335 298062 311344
rect 298008 307760 298060 307766
rect 298008 307702 298060 307708
rect 298020 306649 298048 307702
rect 298006 306640 298062 306649
rect 298006 306575 298062 306584
rect 298008 306332 298060 306338
rect 298008 306274 298060 306280
rect 298020 305289 298048 306274
rect 298006 305280 298062 305289
rect 298006 305215 298062 305224
rect 298572 303929 298600 334698
rect 298744 331696 298796 331702
rect 298744 331638 298796 331644
rect 298650 308680 298706 308689
rect 298650 308615 298706 308624
rect 298558 303920 298614 303929
rect 298558 303855 298614 303864
rect 298008 303544 298060 303550
rect 298008 303486 298060 303492
rect 298020 302569 298048 303486
rect 298006 302560 298062 302569
rect 298006 302495 298062 302504
rect 297822 299160 297878 299169
rect 297822 299095 297878 299104
rect 297744 296686 297864 296714
rect 297730 296440 297786 296449
rect 297730 296375 297786 296384
rect 297744 287178 297772 296375
rect 297836 295186 297864 296686
rect 297824 295180 297876 295186
rect 297824 295122 297876 295128
rect 297822 295080 297878 295089
rect 297822 295015 297878 295024
rect 297836 287434 297864 295015
rect 298008 292528 298060 292534
rect 298008 292470 298060 292476
rect 298020 291689 298048 292470
rect 298006 291680 298062 291689
rect 298006 291615 298062 291624
rect 297914 290320 297970 290329
rect 297914 290255 297970 290264
rect 297928 287450 297956 290255
rect 298008 289672 298060 289678
rect 298008 289614 298060 289620
rect 298020 288969 298048 289614
rect 298006 288960 298062 288969
rect 298006 288895 298062 288904
rect 298008 288380 298060 288386
rect 298008 288322 298060 288328
rect 298020 287609 298048 288322
rect 298006 287600 298062 287609
rect 298006 287535 298062 287544
rect 297824 287428 297876 287434
rect 297928 287422 298048 287450
rect 297824 287370 297876 287376
rect 297744 287150 297956 287178
rect 297824 287088 297876 287094
rect 297824 287030 297876 287036
rect 297836 285938 297864 287030
rect 297824 285932 297876 285938
rect 297824 285874 297876 285880
rect 297928 285818 297956 287150
rect 297744 285790 297956 285818
rect 297638 284200 297694 284209
rect 297638 284135 297694 284144
rect 297744 280634 297772 285790
rect 297824 285728 297876 285734
rect 297824 285670 297876 285676
rect 297732 280628 297784 280634
rect 297732 280570 297784 280576
rect 297548 273964 297600 273970
rect 297548 273906 297600 273912
rect 297640 273284 297692 273290
rect 297640 273226 297692 273232
rect 297364 221536 297416 221542
rect 297364 221478 297416 221484
rect 297272 220176 297324 220182
rect 297272 220118 297324 220124
rect 297284 109993 297312 220118
rect 297270 109984 297326 109993
rect 297270 109919 297326 109928
rect 297376 104009 297404 221478
rect 297454 218240 297510 218249
rect 297454 218175 297510 218184
rect 297362 104000 297418 104009
rect 297362 103935 297418 103944
rect 297468 99521 297496 218175
rect 297548 193180 297600 193186
rect 297548 193122 297600 193128
rect 297560 192273 297588 193122
rect 297546 192264 297602 192273
rect 297546 192199 297602 192208
rect 297548 190460 297600 190466
rect 297548 190402 297600 190408
rect 297560 189281 297588 190402
rect 297546 189272 297602 189281
rect 297546 189207 297602 189216
rect 297546 142896 297602 142905
rect 297546 142831 297602 142840
rect 297560 142186 297588 142831
rect 297548 142180 297600 142186
rect 297548 142122 297600 142128
rect 297652 101017 297680 273226
rect 297730 216200 297786 216209
rect 297730 216135 297786 216144
rect 297744 215354 297772 216135
rect 297732 215348 297784 215354
rect 297732 215290 297784 215296
rect 297730 214704 297786 214713
rect 297730 214639 297786 214648
rect 297744 213994 297772 214639
rect 297732 213988 297784 213994
rect 297732 213930 297784 213936
rect 297730 213208 297786 213217
rect 297730 213143 297786 213152
rect 297744 212566 297772 213143
rect 297732 212560 297784 212566
rect 297732 212502 297784 212508
rect 297730 211712 297786 211721
rect 297730 211647 297786 211656
rect 297744 211206 297772 211647
rect 297732 211200 297784 211206
rect 297732 211142 297784 211148
rect 297730 210216 297786 210225
rect 297730 210151 297786 210160
rect 297744 209846 297772 210151
rect 297732 209840 297784 209846
rect 297732 209782 297784 209788
rect 297730 208720 297786 208729
rect 297730 208655 297786 208664
rect 297744 208418 297772 208655
rect 297732 208412 297784 208418
rect 297732 208354 297784 208360
rect 297730 207224 297786 207233
rect 297730 207159 297786 207168
rect 297744 207058 297772 207159
rect 297732 207052 297784 207058
rect 297732 206994 297784 207000
rect 297730 205728 297786 205737
rect 297730 205663 297732 205672
rect 297784 205663 297786 205672
rect 297732 205634 297784 205640
rect 297730 201240 297786 201249
rect 297730 201175 297786 201184
rect 297744 200190 297772 201175
rect 297732 200184 297784 200190
rect 297732 200126 297784 200132
rect 297730 199744 297786 199753
rect 297730 199679 297786 199688
rect 297744 198762 297772 199679
rect 297732 198756 297784 198762
rect 297732 198698 297784 198704
rect 297730 198248 297786 198257
rect 297730 198183 297786 198192
rect 297744 197402 297772 198183
rect 297732 197396 297784 197402
rect 297732 197338 297784 197344
rect 297730 196752 297786 196761
rect 297730 196687 297786 196696
rect 297744 196042 297772 196687
rect 297732 196036 297784 196042
rect 297732 195978 297784 195984
rect 297730 195256 297786 195265
rect 297730 195191 297786 195200
rect 297744 194614 297772 195191
rect 297732 194608 297784 194614
rect 297732 194550 297784 194556
rect 297730 193760 297786 193769
rect 297730 193695 297786 193704
rect 297744 193254 297772 193695
rect 297732 193248 297784 193254
rect 297732 193190 297784 193196
rect 297730 190768 297786 190777
rect 297730 190703 297786 190712
rect 297744 190534 297772 190703
rect 297732 190528 297784 190534
rect 297732 190470 297784 190476
rect 297732 189032 297784 189038
rect 297732 188974 297784 188980
rect 297744 187785 297772 188974
rect 297730 187776 297786 187785
rect 297730 187711 297786 187720
rect 297732 186312 297784 186318
rect 297730 186280 297732 186289
rect 297784 186280 297786 186289
rect 297730 186215 297786 186224
rect 297732 184884 297784 184890
rect 297732 184826 297784 184832
rect 297744 184793 297772 184826
rect 297730 184784 297786 184793
rect 297730 184719 297786 184728
rect 297732 183524 297784 183530
rect 297732 183466 297784 183472
rect 297744 183297 297772 183466
rect 297730 183288 297786 183297
rect 297730 183223 297786 183232
rect 297732 182164 297784 182170
rect 297732 182106 297784 182112
rect 297744 181801 297772 182106
rect 297730 181792 297786 181801
rect 297730 181727 297786 181736
rect 297732 180804 297784 180810
rect 297732 180746 297784 180752
rect 297744 180305 297772 180746
rect 297730 180296 297786 180305
rect 297730 180231 297786 180240
rect 297732 179376 297784 179382
rect 297732 179318 297784 179324
rect 297744 178809 297772 179318
rect 297730 178800 297786 178809
rect 297730 178735 297786 178744
rect 297732 178016 297784 178022
rect 297732 177958 297784 177964
rect 297744 177313 297772 177958
rect 297730 177304 297786 177313
rect 297730 177239 297786 177248
rect 297732 176656 297784 176662
rect 297732 176598 297784 176604
rect 297744 175817 297772 176598
rect 297730 175808 297786 175817
rect 297730 175743 297786 175752
rect 297732 175228 297784 175234
rect 297732 175170 297784 175176
rect 297744 174321 297772 175170
rect 297730 174312 297786 174321
rect 297730 174247 297786 174256
rect 297732 173188 297784 173194
rect 297732 173130 297784 173136
rect 297744 172825 297772 173130
rect 297730 172816 297786 172825
rect 297730 172751 297786 172760
rect 297730 171320 297786 171329
rect 297730 171255 297786 171264
rect 297744 171154 297772 171255
rect 297732 171148 297784 171154
rect 297732 171090 297784 171096
rect 297730 169824 297786 169833
rect 297730 169759 297732 169768
rect 297784 169759 297786 169768
rect 297732 169730 297784 169736
rect 297730 168328 297786 168337
rect 297730 168263 297786 168272
rect 297744 167074 297772 168263
rect 297732 167068 297784 167074
rect 297732 167010 297784 167016
rect 297730 165336 297786 165345
rect 297730 165271 297786 165280
rect 297744 164286 297772 165271
rect 297732 164280 297784 164286
rect 297732 164222 297784 164228
rect 297730 163840 297786 163849
rect 297730 163775 297786 163784
rect 297744 162926 297772 163775
rect 297732 162920 297784 162926
rect 297732 162862 297784 162868
rect 297730 162344 297786 162353
rect 297730 162279 297786 162288
rect 297744 161498 297772 162279
rect 297732 161492 297784 161498
rect 297732 161434 297784 161440
rect 297730 160848 297786 160857
rect 297730 160783 297786 160792
rect 297744 160138 297772 160783
rect 297732 160132 297784 160138
rect 297732 160074 297784 160080
rect 297730 159352 297786 159361
rect 297730 159287 297786 159296
rect 297744 158778 297772 159287
rect 297732 158772 297784 158778
rect 297732 158714 297784 158720
rect 297730 156360 297786 156369
rect 297730 156295 297786 156304
rect 297744 155990 297772 156295
rect 297732 155984 297784 155990
rect 297732 155926 297784 155932
rect 297730 154864 297786 154873
rect 297730 154799 297786 154808
rect 297744 154630 297772 154799
rect 297732 154624 297784 154630
rect 297732 154566 297784 154572
rect 297730 153368 297786 153377
rect 297730 153303 297786 153312
rect 297744 153270 297772 153303
rect 297732 153264 297784 153270
rect 297732 153206 297784 153212
rect 297730 151872 297786 151881
rect 297730 151807 297732 151816
rect 297784 151807 297786 151816
rect 297732 151778 297784 151784
rect 297730 150376 297786 150385
rect 297730 150311 297786 150320
rect 297744 149122 297772 150311
rect 297732 149116 297784 149122
rect 297732 149058 297784 149064
rect 297730 147384 297786 147393
rect 297730 147319 297786 147328
rect 297744 146334 297772 147319
rect 297732 146328 297784 146334
rect 297732 146270 297784 146276
rect 297730 145888 297786 145897
rect 297730 145823 297786 145832
rect 297744 144974 297772 145823
rect 297732 144968 297784 144974
rect 297732 144910 297784 144916
rect 297730 144392 297786 144401
rect 297730 144327 297786 144336
rect 297744 143614 297772 144327
rect 297732 143608 297784 143614
rect 297732 143550 297784 143556
rect 297732 142112 297784 142118
rect 297732 142054 297784 142060
rect 297744 141409 297772 142054
rect 297730 141400 297786 141409
rect 297730 141335 297786 141344
rect 297732 140752 297784 140758
rect 297732 140694 297784 140700
rect 297744 139913 297772 140694
rect 297730 139904 297786 139913
rect 297730 139839 297786 139848
rect 297732 139392 297784 139398
rect 297732 139334 297784 139340
rect 297744 138417 297772 139334
rect 297730 138408 297786 138417
rect 297730 138343 297786 138352
rect 297732 137964 297784 137970
rect 297732 137906 297784 137912
rect 297744 136921 297772 137906
rect 297730 136912 297786 136921
rect 297730 136847 297786 136856
rect 297732 135244 297784 135250
rect 297732 135186 297784 135192
rect 297744 133929 297772 135186
rect 297730 133920 297786 133929
rect 297730 133855 297786 133864
rect 297732 132456 297784 132462
rect 297730 132424 297732 132433
rect 297784 132424 297786 132433
rect 297730 132359 297786 132368
rect 297732 131096 297784 131102
rect 297732 131038 297784 131044
rect 297744 130937 297772 131038
rect 297730 130928 297786 130937
rect 297730 130863 297786 130872
rect 297732 129736 297784 129742
rect 297732 129678 297784 129684
rect 297744 129441 297772 129678
rect 297730 129432 297786 129441
rect 297730 129367 297786 129376
rect 297732 128308 297784 128314
rect 297732 128250 297784 128256
rect 297744 127945 297772 128250
rect 297730 127936 297786 127945
rect 297730 127871 297786 127880
rect 297732 126948 297784 126954
rect 297732 126890 297784 126896
rect 297744 126449 297772 126890
rect 297730 126440 297786 126449
rect 297730 126375 297786 126384
rect 297732 125588 297784 125594
rect 297732 125530 297784 125536
rect 297744 124953 297772 125530
rect 297730 124944 297786 124953
rect 297730 124879 297786 124888
rect 297732 124160 297784 124166
rect 297732 124102 297784 124108
rect 297744 123457 297772 124102
rect 297730 123448 297786 123457
rect 297730 123383 297786 123392
rect 297732 122800 297784 122806
rect 297732 122742 297784 122748
rect 297744 121961 297772 122742
rect 297730 121952 297786 121961
rect 297730 121887 297786 121896
rect 297732 121440 297784 121446
rect 297732 121382 297784 121388
rect 297744 120465 297772 121382
rect 297730 120456 297786 120465
rect 297730 120391 297786 120400
rect 297732 120080 297784 120086
rect 297732 120022 297784 120028
rect 297744 118969 297772 120022
rect 297730 118960 297786 118969
rect 297730 118895 297786 118904
rect 297732 117292 297784 117298
rect 297732 117234 297784 117240
rect 297744 115977 297772 117234
rect 297730 115968 297786 115977
rect 297730 115903 297786 115912
rect 297732 114504 297784 114510
rect 297730 114472 297732 114481
rect 297784 114472 297786 114481
rect 297730 114407 297786 114416
rect 297732 113144 297784 113150
rect 297732 113086 297784 113092
rect 297744 112985 297772 113086
rect 297730 112976 297786 112985
rect 297730 112911 297786 112920
rect 297638 101008 297694 101017
rect 297638 100943 297694 100952
rect 297454 99512 297510 99521
rect 297454 99447 297510 99456
rect 297836 96529 297864 285670
rect 297916 285660 297968 285666
rect 297916 285602 297968 285608
rect 297928 285569 297956 285602
rect 297914 285560 297970 285569
rect 297914 285495 297970 285504
rect 297916 276072 297968 276078
rect 297916 276014 297968 276020
rect 297928 107001 297956 276014
rect 297914 106992 297970 107001
rect 297914 106927 297970 106936
rect 297822 96520 297878 96529
rect 297822 96455 297878 96464
rect 297086 92032 297142 92041
rect 297086 91967 297142 91976
rect 298020 90545 298048 287422
rect 298664 278050 298692 308615
rect 298652 278044 298704 278050
rect 298652 277986 298704 277992
rect 298756 273290 298784 331638
rect 298836 331492 298888 331498
rect 298836 331434 298888 331440
rect 298848 276078 298876 331434
rect 298928 331356 298980 331362
rect 298928 331298 298980 331304
rect 298940 279954 298968 331298
rect 299032 281353 299060 348366
rect 299492 337550 299520 494634
rect 299572 454028 299624 454034
rect 299572 453970 299624 453976
rect 299480 337544 299532 337550
rect 299480 337486 299532 337492
rect 299204 330132 299256 330138
rect 299204 330074 299256 330080
rect 299112 329996 299164 330002
rect 299112 329938 299164 329944
rect 299018 281344 299074 281353
rect 299018 281279 299074 281288
rect 298928 279948 298980 279954
rect 298928 279890 298980 279896
rect 298836 276072 298888 276078
rect 298836 276014 298888 276020
rect 298744 273284 298796 273290
rect 298744 273226 298796 273232
rect 298928 221604 298980 221610
rect 298928 221546 298980 221552
rect 298836 220244 298888 220250
rect 298836 220186 298888 220192
rect 298848 98025 298876 220186
rect 298834 98016 298890 98025
rect 298834 97951 298890 97960
rect 298940 93537 298968 221546
rect 299020 220312 299072 220318
rect 299020 220254 299072 220260
rect 298926 93528 298982 93537
rect 298926 93463 298982 93472
rect 298006 90536 298062 90545
rect 298006 90471 298062 90480
rect 296812 90364 296864 90370
rect 296812 90306 296864 90312
rect 296824 86057 296852 90306
rect 299032 89049 299060 220254
rect 299124 111489 299152 329938
rect 299110 111480 299166 111489
rect 299110 111415 299166 111424
rect 299216 108497 299244 330074
rect 299296 330064 299348 330070
rect 299296 330006 299348 330012
rect 299202 108488 299258 108497
rect 299202 108423 299258 108432
rect 299308 105505 299336 330006
rect 299388 329928 299440 329934
rect 299388 329870 299440 329876
rect 299294 105496 299350 105505
rect 299294 105431 299350 105440
rect 299400 95033 299428 329870
rect 299584 297809 299612 453970
rect 299676 362234 299704 500126
rect 299848 496868 299900 496874
rect 299848 496810 299900 496816
rect 299664 362228 299716 362234
rect 299664 362170 299716 362176
rect 299662 322280 299718 322289
rect 299662 322215 299718 322224
rect 299570 297800 299626 297809
rect 299570 297735 299626 297744
rect 299570 282840 299626 282849
rect 299570 282775 299626 282784
rect 299478 281480 299534 281489
rect 299478 281415 299534 281424
rect 299492 222154 299520 281415
rect 299584 275330 299612 282775
rect 299572 275324 299624 275330
rect 299572 275266 299624 275272
rect 299676 271862 299704 322215
rect 299756 295180 299808 295186
rect 299756 295122 299808 295128
rect 299664 271856 299716 271862
rect 299664 271798 299716 271804
rect 299768 223106 299796 295122
rect 299860 280022 299888 496810
rect 300412 494698 300440 500126
rect 300400 494692 300452 494698
rect 300400 494634 300452 494640
rect 300964 454034 300992 500126
rect 301884 497758 301912 500126
rect 301872 497752 301924 497758
rect 301872 497694 301924 497700
rect 302332 492652 302384 492658
rect 302332 492594 302384 492600
rect 300952 454028 301004 454034
rect 300952 453970 301004 453976
rect 301504 371272 301556 371278
rect 301504 371214 301556 371220
rect 301516 333198 301544 371214
rect 301504 333192 301556 333198
rect 301504 333134 301556 333140
rect 300674 331664 300730 331673
rect 300674 331599 300730 331608
rect 300688 329868 300716 331599
rect 301964 331288 302016 331294
rect 301964 331230 302016 331236
rect 301976 329868 302004 331230
rect 302344 330018 302372 492594
rect 302436 331906 302464 500126
rect 303678 499882 303706 500140
rect 303632 499854 303706 499882
rect 303816 500126 304428 500154
rect 303632 331906 303660 499854
rect 303816 341630 303844 500126
rect 305150 499882 305178 500140
rect 305104 499854 305178 499882
rect 305564 500126 305900 500154
rect 306392 500126 306636 500154
rect 306760 500126 307372 500154
rect 307864 500126 308108 500154
rect 308508 500126 308844 500154
rect 309152 500126 309580 500154
rect 309704 500126 310316 500154
rect 310532 500126 311052 500154
rect 311176 500126 311788 500154
rect 312004 500126 312524 500154
rect 312924 500126 313260 500154
rect 313384 500126 313996 500154
rect 303804 341624 303856 341630
rect 303804 341566 303856 341572
rect 305104 332178 305132 499854
rect 305564 496874 305592 500126
rect 305552 496868 305604 496874
rect 305552 496810 305604 496816
rect 305092 332172 305144 332178
rect 305092 332114 305144 332120
rect 306392 332110 306420 500126
rect 306760 489914 306788 500126
rect 307760 494692 307812 494698
rect 307760 494634 307812 494640
rect 306484 489886 306788 489914
rect 306484 333402 306512 489886
rect 307772 348430 307800 494634
rect 307864 355366 307892 500126
rect 308508 494698 308536 500126
rect 308496 494692 308548 494698
rect 308496 494634 308548 494640
rect 307852 355360 307904 355366
rect 307852 355302 307904 355308
rect 307760 348424 307812 348430
rect 307760 348366 307812 348372
rect 306472 333396 306524 333402
rect 306472 333338 306524 333344
rect 306472 333192 306524 333198
rect 306472 333134 306524 333140
rect 306380 332104 306432 332110
rect 306380 332046 306432 332052
rect 302424 331900 302476 331906
rect 302424 331842 302476 331848
rect 303620 331900 303672 331906
rect 303620 331842 303672 331848
rect 305182 331256 305238 331265
rect 305182 331191 305238 331200
rect 302344 329990 302832 330018
rect 302804 329882 302832 329990
rect 302804 329854 303278 329882
rect 305196 329868 305224 331191
rect 306484 329868 306512 333134
rect 309152 332042 309180 500126
rect 309704 489914 309732 500126
rect 309244 489886 309732 489914
rect 309140 332036 309192 332042
rect 309140 331978 309192 331984
rect 309244 331974 309272 489886
rect 310532 334694 310560 500126
rect 311176 489914 311204 500126
rect 311900 494352 311952 494358
rect 311900 494294 311952 494300
rect 310624 489886 311204 489914
rect 310624 480962 310652 489886
rect 310612 480956 310664 480962
rect 310612 480898 310664 480904
rect 311912 334762 311940 494294
rect 312004 344418 312032 500126
rect 312924 494358 312952 500126
rect 312912 494352 312964 494358
rect 312912 494294 312964 494300
rect 313384 460222 313412 500126
rect 314718 499882 314746 500140
rect 314672 499854 314746 499882
rect 315132 500126 315468 500154
rect 316052 500126 316204 500154
rect 316604 500126 316940 500154
rect 317432 500126 317676 500154
rect 314672 497554 314700 499854
rect 315132 497894 315160 500126
rect 316052 497962 316080 500126
rect 316040 497956 316092 497962
rect 316040 497898 316092 497904
rect 315120 497888 315172 497894
rect 315120 497830 315172 497836
rect 316604 497690 316632 500126
rect 316592 497684 316644 497690
rect 316592 497626 316644 497632
rect 317432 497622 317460 500126
rect 317420 497616 317472 497622
rect 317420 497558 317472 497564
rect 314660 497548 314712 497554
rect 314660 497490 314712 497496
rect 313372 460216 313424 460222
rect 313372 460158 313424 460164
rect 313924 389224 313976 389230
rect 313924 389166 313976 389172
rect 311992 344412 312044 344418
rect 311992 344354 312044 344360
rect 311992 341692 312044 341698
rect 311992 341634 312044 341640
rect 311900 334756 311952 334762
rect 311900 334698 311952 334704
rect 310520 334688 310572 334694
rect 310520 334630 310572 334636
rect 310334 332208 310390 332217
rect 310334 332143 310390 332152
rect 309232 331968 309284 331974
rect 309232 331910 309284 331916
rect 309048 331764 309100 331770
rect 309048 331706 309100 331712
rect 307760 331356 307812 331362
rect 307760 331298 307812 331304
rect 307772 329868 307800 331298
rect 309060 329868 309088 331706
rect 310348 329868 310376 332143
rect 312004 329882 312032 341634
rect 313936 335442 313964 389166
rect 314660 362228 314712 362234
rect 314660 362170 314712 362176
rect 313924 335436 313976 335442
rect 313924 335378 313976 335384
rect 313556 331628 313608 331634
rect 313556 331570 313608 331576
rect 312004 329854 312294 329882
rect 313568 329868 313596 331570
rect 314672 329882 314700 362170
rect 318904 338842 318932 505514
rect 318996 344350 319024 506466
rect 319088 345710 319116 507826
rect 319180 351218 319208 509206
rect 320180 509186 320232 509192
rect 319350 508328 319406 508337
rect 319350 508263 319352 508272
rect 319404 508263 319406 508272
rect 319352 508234 319404 508240
rect 320192 508133 320220 509186
rect 320178 508124 320234 508133
rect 320178 508059 320234 508068
rect 320364 507816 320416 507822
rect 320364 507758 320416 507764
rect 320088 507680 320140 507686
rect 320088 507622 320140 507628
rect 320100 506773 320128 507622
rect 320376 507453 320404 507758
rect 320362 507444 320418 507453
rect 320284 507402 320362 507430
rect 320086 506764 320142 506773
rect 320086 506699 320142 506708
rect 320100 506530 320128 506699
rect 320088 506524 320140 506530
rect 320088 506466 320140 506472
rect 320180 506456 320232 506462
rect 320180 506398 320232 506404
rect 319352 505776 319404 505782
rect 319352 505718 319404 505724
rect 319364 505617 319392 505718
rect 319350 505608 319406 505617
rect 319350 505543 319352 505552
rect 319404 505543 319406 505552
rect 319352 505514 319404 505520
rect 320192 505413 320220 506398
rect 320178 505404 320234 505413
rect 320178 505339 320234 505348
rect 320192 505170 320220 505339
rect 320180 505164 320232 505170
rect 320180 505106 320232 505112
rect 320088 505028 320140 505034
rect 320088 504970 320140 504976
rect 320100 504733 320128 504970
rect 320086 504724 320142 504733
rect 320086 504659 320142 504668
rect 319350 504248 319406 504257
rect 319350 504183 319406 504192
rect 319364 489914 319392 504183
rect 320180 503668 320232 503674
rect 320180 503610 320232 503616
rect 319272 489886 319392 489914
rect 319168 351212 319220 351218
rect 319168 351154 319220 351160
rect 319076 345704 319128 345710
rect 319076 345646 319128 345652
rect 318984 344344 319036 344350
rect 318984 344286 319036 344292
rect 318892 338836 318944 338842
rect 318892 338778 318944 338784
rect 319272 337414 319300 489886
rect 319352 337544 319404 337550
rect 319352 337486 319404 337492
rect 319260 337408 319312 337414
rect 319260 337350 319312 337356
rect 318064 335436 318116 335442
rect 318064 335378 318116 335384
rect 316130 331392 316186 331401
rect 316130 331327 316186 331336
rect 314672 329854 314870 329882
rect 316144 329868 316172 331327
rect 318076 329868 318104 335378
rect 319364 329868 319392 337486
rect 320192 333266 320220 503610
rect 320284 499574 320312 507402
rect 320362 507379 320418 507388
rect 320284 499546 320404 499574
rect 320376 487830 320404 499546
rect 320468 494766 320496 509487
rect 320546 508056 320602 508065
rect 320546 507991 320602 508000
rect 320560 496194 320588 507991
rect 320652 500274 320680 510818
rect 320732 505164 320784 505170
rect 320732 505106 320784 505112
rect 320640 500268 320692 500274
rect 320640 500210 320692 500216
rect 320548 496188 320600 496194
rect 320548 496130 320600 496136
rect 320744 496126 320772 505106
rect 320732 496120 320784 496126
rect 320732 496062 320784 496068
rect 320456 494760 320508 494766
rect 320456 494702 320508 494708
rect 320364 487824 320416 487830
rect 320364 487766 320416 487772
rect 320836 365702 320864 640358
rect 320928 565049 320956 700402
rect 321100 642320 321152 642326
rect 321100 642262 321152 642268
rect 321008 642116 321060 642122
rect 321008 642058 321060 642064
rect 320914 565040 320970 565049
rect 320914 564975 320970 564984
rect 321020 555393 321048 642058
rect 321112 561134 321140 642262
rect 323676 642252 323728 642258
rect 323676 642194 323728 642200
rect 322388 640484 322440 640490
rect 322388 640426 322440 640432
rect 322204 639124 322256 639130
rect 322204 639066 322256 639072
rect 321100 561128 321152 561134
rect 321100 561070 321152 561076
rect 321006 555384 321062 555393
rect 321006 555319 321062 555328
rect 322216 552770 322244 639066
rect 322296 638988 322348 638994
rect 322296 638930 322348 638936
rect 322308 552906 322336 638930
rect 322400 578202 322428 640426
rect 323584 640348 323636 640354
rect 323584 640290 323636 640296
rect 322480 639396 322532 639402
rect 322480 639338 322532 639344
rect 322492 585818 322520 639338
rect 322480 585812 322532 585818
rect 322480 585754 322532 585760
rect 322388 578196 322440 578202
rect 322388 578138 322440 578144
rect 322296 552900 322348 552906
rect 322296 552842 322348 552848
rect 322204 552764 322256 552770
rect 322204 552706 322256 552712
rect 322204 549908 322256 549914
rect 322204 549850 322256 549856
rect 322216 535401 322244 549850
rect 322296 548616 322348 548622
rect 322296 548558 322348 548564
rect 322202 535392 322258 535401
rect 322202 535327 322258 535336
rect 321652 532704 321704 532710
rect 321652 532646 321704 532652
rect 321664 532273 321692 532646
rect 322202 532400 322258 532409
rect 322202 532335 322258 532344
rect 321650 532264 321706 532273
rect 321650 532199 321706 532208
rect 321560 527264 321612 527270
rect 321560 527206 321612 527212
rect 321572 527105 321600 527206
rect 321558 527096 321614 527105
rect 321558 527031 321614 527040
rect 322020 522980 322072 522986
rect 322020 522922 322072 522928
rect 322032 521937 322060 522922
rect 322018 521928 322074 521937
rect 322018 521863 322074 521872
rect 322020 521620 322072 521626
rect 322020 521562 322072 521568
rect 322032 520577 322060 521562
rect 322018 520568 322074 520577
rect 322018 520503 322074 520512
rect 321558 519344 321614 519353
rect 321558 519279 321560 519288
rect 321612 519279 321614 519288
rect 321560 519250 321612 519256
rect 321836 518900 321888 518906
rect 321836 518842 321888 518848
rect 321848 517857 321876 518842
rect 321834 517848 321890 517857
rect 321834 517783 321890 517792
rect 321560 517472 321612 517478
rect 321558 517440 321560 517449
rect 321612 517440 321614 517449
rect 321558 517375 321614 517384
rect 321836 516112 321888 516118
rect 321836 516054 321888 516060
rect 321848 515409 321876 516054
rect 321834 515400 321890 515409
rect 321834 515335 321890 515344
rect 321650 514176 321706 514185
rect 321650 514111 321706 514120
rect 322110 514176 322166 514185
rect 322110 514111 322166 514120
rect 320914 512136 320970 512145
rect 320914 512071 320970 512080
rect 320824 365696 320876 365702
rect 320824 365638 320876 365644
rect 320272 341624 320324 341630
rect 320272 341566 320324 341572
rect 320180 333260 320232 333266
rect 320180 333202 320232 333208
rect 320284 329882 320312 341566
rect 320928 340105 320956 512071
rect 321558 511320 321614 511329
rect 321558 511255 321560 511264
rect 321612 511255 321614 511264
rect 321560 511226 321612 511232
rect 320914 340096 320970 340105
rect 320914 340031 320970 340040
rect 321572 334665 321600 511226
rect 321664 500342 321692 514111
rect 322124 514078 322152 514111
rect 322112 514072 322164 514078
rect 322112 514014 322164 514020
rect 321742 512680 321798 512689
rect 321742 512615 321798 512624
rect 322110 512680 322166 512689
rect 322110 512615 322112 512624
rect 321756 500410 321784 512615
rect 322164 512615 322166 512624
rect 322112 512586 322164 512592
rect 321744 500404 321796 500410
rect 321744 500346 321796 500352
rect 321652 500336 321704 500342
rect 321652 500278 321704 500284
rect 322216 500274 322244 532335
rect 322308 528465 322336 548558
rect 322478 536208 322534 536217
rect 322478 536143 322534 536152
rect 322388 536104 322440 536110
rect 322388 536046 322440 536052
rect 322400 534041 322428 536046
rect 322492 534750 322520 536143
rect 322480 534744 322532 534750
rect 322480 534686 322532 534692
rect 322478 534440 322534 534449
rect 322478 534375 322534 534384
rect 322492 534138 322520 534375
rect 322480 534132 322532 534138
rect 322480 534074 322532 534080
rect 322386 534032 322442 534041
rect 322386 533967 322442 533976
rect 322848 533452 322900 533458
rect 322848 533394 322900 533400
rect 322860 533361 322888 533394
rect 322846 533352 322902 533361
rect 322846 533287 322902 533296
rect 322480 531208 322532 531214
rect 322478 531176 322480 531185
rect 322532 531176 322534 531185
rect 322478 531111 322534 531120
rect 322386 530224 322442 530233
rect 322386 530159 322442 530168
rect 322400 529990 322428 530159
rect 322388 529984 322440 529990
rect 322388 529926 322440 529932
rect 322480 529916 322532 529922
rect 322480 529858 322532 529864
rect 322492 529825 322520 529858
rect 322478 529816 322534 529825
rect 322478 529751 322534 529760
rect 322860 529242 322888 533287
rect 322848 529236 322900 529242
rect 322848 529178 322900 529184
rect 322754 528864 322810 528873
rect 322754 528799 322810 528808
rect 322480 528556 322532 528562
rect 322480 528498 322532 528504
rect 322294 528456 322350 528465
rect 322294 528391 322350 528400
rect 322492 528193 322520 528498
rect 322478 528184 322534 528193
rect 322478 528119 322534 528128
rect 322480 527128 322532 527134
rect 322480 527070 322532 527076
rect 322492 526833 322520 527070
rect 322478 526824 322534 526833
rect 322478 526759 322534 526768
rect 322480 525768 322532 525774
rect 322478 525736 322480 525745
rect 322532 525736 322534 525745
rect 322478 525671 322534 525680
rect 322768 525094 322796 528799
rect 322756 525088 322808 525094
rect 322756 525030 322808 525036
rect 322570 524648 322626 524657
rect 322570 524583 322626 524592
rect 322294 524512 322350 524521
rect 322294 524447 322350 524456
rect 322204 500268 322256 500274
rect 322204 500210 322256 500216
rect 322308 499390 322336 524447
rect 322478 523424 322534 523433
rect 322478 523359 322534 523368
rect 322386 523152 322442 523161
rect 322386 523087 322442 523096
rect 322400 516798 322428 523087
rect 322492 523054 322520 523359
rect 322480 523048 322532 523054
rect 322480 522990 322532 522996
rect 322478 522064 322534 522073
rect 322478 521999 322534 522008
rect 322492 521694 322520 521999
rect 322480 521688 322532 521694
rect 322480 521630 322532 521636
rect 322478 520704 322534 520713
rect 322478 520639 322534 520648
rect 322492 520334 322520 520639
rect 322480 520328 322532 520334
rect 322480 520270 322532 520276
rect 322478 517984 322534 517993
rect 322478 517919 322534 517928
rect 322492 517614 322520 517919
rect 322480 517608 322532 517614
rect 322480 517550 322532 517556
rect 322388 516792 322440 516798
rect 322388 516734 322440 516740
rect 322388 516384 322440 516390
rect 322386 516352 322388 516361
rect 322440 516352 322442 516361
rect 322386 516287 322442 516296
rect 322478 513496 322534 513505
rect 322478 513431 322534 513440
rect 322492 513398 322520 513431
rect 322480 513392 322532 513398
rect 322480 513334 322532 513340
rect 322584 509234 322612 524583
rect 322848 519580 322900 519586
rect 322848 519522 322900 519528
rect 322860 519217 322888 519522
rect 322846 519208 322902 519217
rect 322846 519143 322902 519152
rect 322940 516384 322992 516390
rect 322940 516326 322992 516332
rect 322846 515536 322902 515545
rect 322846 515471 322902 515480
rect 322860 515438 322888 515471
rect 322848 515432 322900 515438
rect 322848 515374 322900 515380
rect 322492 509206 322612 509234
rect 322388 504212 322440 504218
rect 322388 504154 322440 504160
rect 322400 504121 322428 504154
rect 322386 504112 322442 504121
rect 322386 504047 322442 504056
rect 322388 503600 322440 503606
rect 322388 503542 322440 503548
rect 322400 503441 322428 503542
rect 322386 503432 322442 503441
rect 322386 503367 322442 503376
rect 322386 502480 322442 502489
rect 322386 502415 322442 502424
rect 322400 502382 322428 502415
rect 322388 502376 322440 502382
rect 322388 502318 322440 502324
rect 322296 499384 322348 499390
rect 322296 499326 322348 499332
rect 322492 498846 322520 509206
rect 322480 498840 322532 498846
rect 322480 498782 322532 498788
rect 321558 334656 321614 334665
rect 321558 334591 321614 334600
rect 322952 331809 322980 516326
rect 323596 419490 323624 640290
rect 323688 574802 323716 642194
rect 329196 642184 329248 642190
rect 329196 642126 329248 642132
rect 325056 641980 325108 641986
rect 325056 641922 325108 641928
rect 324964 598188 325016 598194
rect 324964 598130 325016 598136
rect 324228 594176 324280 594182
rect 324228 594118 324280 594124
rect 323676 574796 323728 574802
rect 323676 574738 323728 574744
rect 323676 543040 323728 543046
rect 323676 542982 323728 542988
rect 323688 527270 323716 542982
rect 323768 532772 323820 532778
rect 323768 532714 323820 532720
rect 323676 527264 323728 527270
rect 323676 527206 323728 527212
rect 323676 519308 323728 519314
rect 323676 519250 323728 519256
rect 323688 498914 323716 519250
rect 323780 517478 323808 532714
rect 324240 519586 324268 594118
rect 324228 519580 324280 519586
rect 324228 519522 324280 519528
rect 323768 517472 323820 517478
rect 323768 517414 323820 517420
rect 324228 515432 324280 515438
rect 324228 515374 324280 515380
rect 324240 509930 324268 515374
rect 324228 509924 324280 509930
rect 324228 509866 324280 509872
rect 323676 498908 323728 498914
rect 323676 498850 323728 498856
rect 324976 498642 325004 598130
rect 325068 552702 325096 641922
rect 327724 639736 327776 639742
rect 327724 639678 327776 639684
rect 327736 596970 327764 639678
rect 327724 596964 327776 596970
rect 327724 596906 327776 596912
rect 327724 596828 327776 596834
rect 327724 596770 327776 596776
rect 329104 596828 329156 596834
rect 329104 596770 329156 596776
rect 325516 591388 325568 591394
rect 325516 591330 325568 591336
rect 325056 552696 325108 552702
rect 325056 552638 325108 552644
rect 325056 549296 325108 549302
rect 325056 549238 325108 549244
rect 325068 516390 325096 549238
rect 325056 516384 325108 516390
rect 325056 516326 325108 516332
rect 325528 505782 325556 591330
rect 326988 549364 327040 549370
rect 326988 549306 327040 549312
rect 325608 537532 325660 537538
rect 325608 537474 325660 537480
rect 325516 505776 325568 505782
rect 325516 505718 325568 505724
rect 325620 503674 325648 537474
rect 327000 518945 327028 549306
rect 325698 518936 325754 518945
rect 325698 518871 325700 518880
rect 325752 518871 325754 518880
rect 326986 518936 327042 518945
rect 326986 518871 327042 518880
rect 325700 518842 325752 518848
rect 326344 517540 326396 517546
rect 326344 517482 326396 517488
rect 326356 504218 326384 517482
rect 327736 505102 327764 596770
rect 327816 594108 327868 594114
rect 327816 594050 327868 594056
rect 327828 532642 327856 594050
rect 327906 541104 327962 541113
rect 327906 541039 327962 541048
rect 327816 532636 327868 532642
rect 327816 532578 327868 532584
rect 327920 510882 327948 541039
rect 329116 537538 329144 596770
rect 329104 537532 329156 537538
rect 329104 537474 329156 537480
rect 328368 533384 328420 533390
rect 328368 533326 328420 533332
rect 328380 531214 328408 533326
rect 328368 531208 328420 531214
rect 328368 531150 328420 531156
rect 329208 513262 329236 642126
rect 331232 594114 331260 702986
rect 348804 702434 348832 703520
rect 347792 702406 348832 702434
rect 337384 697604 337436 697610
rect 337384 697546 337436 697552
rect 331864 642048 331916 642054
rect 331864 641990 331916 641996
rect 333244 642048 333296 642054
rect 333244 641990 333296 641996
rect 331220 594108 331272 594114
rect 331220 594050 331272 594056
rect 329288 587172 329340 587178
rect 329288 587114 329340 587120
rect 329300 515438 329328 587114
rect 330484 540252 330536 540258
rect 330484 540194 330536 540200
rect 330496 539578 330524 540194
rect 330484 539572 330536 539578
rect 330484 539514 330536 539520
rect 330484 534744 330536 534750
rect 330484 534686 330536 534692
rect 330496 530641 330524 534686
rect 330482 530632 330538 530641
rect 330482 530567 330538 530576
rect 331876 527066 331904 641990
rect 333256 599350 333284 641990
rect 333244 599344 333296 599350
rect 333244 599286 333296 599292
rect 336004 596896 336056 596902
rect 336004 596838 336056 596844
rect 334624 595604 334676 595610
rect 334624 595546 334676 595552
rect 333888 595536 333940 595542
rect 333888 595478 333940 595484
rect 331956 594244 332008 594250
rect 331956 594186 332008 594192
rect 331864 527060 331916 527066
rect 331864 527002 331916 527008
rect 329288 515432 329340 515438
rect 329288 515374 329340 515380
rect 331968 514758 331996 594186
rect 333244 590028 333296 590034
rect 333244 589970 333296 589976
rect 332046 547088 332102 547097
rect 332046 547023 332102 547032
rect 331956 514752 332008 514758
rect 331956 514694 332008 514700
rect 332060 514078 332088 547023
rect 333256 524414 333284 589970
rect 333900 550730 333928 595478
rect 333336 550724 333388 550730
rect 333336 550666 333388 550672
rect 333888 550724 333940 550730
rect 333888 550666 333940 550672
rect 333244 524408 333296 524414
rect 333244 524350 333296 524356
rect 332048 514072 332100 514078
rect 332048 514014 332100 514020
rect 329196 513256 329248 513262
rect 329196 513198 329248 513204
rect 327908 510876 327960 510882
rect 327908 510818 327960 510824
rect 333348 510542 333376 550666
rect 333336 510536 333388 510542
rect 333336 510478 333388 510484
rect 334636 507754 334664 595546
rect 336016 532574 336044 596838
rect 336648 590028 336700 590034
rect 336648 589970 336700 589976
rect 336004 532568 336056 532574
rect 336004 532510 336056 532516
rect 336660 511290 336688 589970
rect 336648 511284 336700 511290
rect 336648 511226 336700 511232
rect 334624 507748 334676 507754
rect 334624 507690 334676 507696
rect 327724 505096 327776 505102
rect 327724 505038 327776 505044
rect 326344 504212 326396 504218
rect 326344 504154 326396 504160
rect 325608 503668 325660 503674
rect 325608 503610 325660 503616
rect 337396 502314 337424 697546
rect 338764 640688 338816 640694
rect 338764 640630 338816 640636
rect 342904 640688 342956 640694
rect 342904 640630 342956 640636
rect 337476 569288 337528 569294
rect 337476 569230 337528 569236
rect 337488 529854 337516 569230
rect 337476 529848 337528 529854
rect 337476 529790 337528 529796
rect 337568 529236 337620 529242
rect 337568 529178 337620 529184
rect 337580 510542 337608 529178
rect 337568 510536 337620 510542
rect 337568 510478 337620 510484
rect 337384 502308 337436 502314
rect 337384 502250 337436 502256
rect 324964 498636 325016 498642
rect 324964 498578 325016 498584
rect 327724 497820 327776 497826
rect 327724 497762 327776 497768
rect 323676 423700 323728 423706
rect 323676 423642 323728 423648
rect 323584 419484 323636 419490
rect 323584 419426 323636 419432
rect 323216 332240 323268 332246
rect 323216 332182 323268 332188
rect 322938 331800 322994 331809
rect 322938 331735 322994 331744
rect 321928 331560 321980 331566
rect 321928 331502 321980 331508
rect 320284 329854 320666 329882
rect 321940 329868 321968 331502
rect 323228 329868 323256 332182
rect 323688 331838 323716 423642
rect 323676 331832 323728 331838
rect 323676 331774 323728 331780
rect 325148 331832 325200 331838
rect 325148 331774 325200 331780
rect 325160 329868 325188 331774
rect 327736 331566 327764 497762
rect 338776 471986 338804 640630
rect 342916 598602 342944 640630
rect 342904 598596 342956 598602
rect 342904 598538 342956 598544
rect 342168 596896 342220 596902
rect 342168 596838 342220 596844
rect 338856 588668 338908 588674
rect 338856 588610 338908 588616
rect 338868 535430 338896 588610
rect 340144 584588 340196 584594
rect 340144 584530 340196 584536
rect 338856 535424 338908 535430
rect 338856 535366 338908 535372
rect 340156 533458 340184 584530
rect 341524 548548 341576 548554
rect 341524 548490 341576 548496
rect 340236 541748 340288 541754
rect 340236 541690 340288 541696
rect 340144 533452 340196 533458
rect 340144 533394 340196 533400
rect 340248 511970 340276 541690
rect 340880 536852 340932 536858
rect 340880 536794 340932 536800
rect 340892 536110 340920 536794
rect 340880 536104 340932 536110
rect 340880 536046 340932 536052
rect 341536 517478 341564 548490
rect 341524 517472 341576 517478
rect 341524 517414 341576 517420
rect 340236 511964 340288 511970
rect 340236 511906 340288 511912
rect 342180 505170 342208 596838
rect 347792 595474 347820 702406
rect 360844 700460 360896 700466
rect 360844 700402 360896 700408
rect 355416 663876 355468 663882
rect 355416 663818 355468 663824
rect 352564 663808 352616 663814
rect 352564 663750 352616 663756
rect 351368 642388 351420 642394
rect 351368 642330 351420 642336
rect 349896 642252 349948 642258
rect 349896 642194 349948 642200
rect 349804 641844 349856 641850
rect 349804 641786 349856 641792
rect 345664 595468 345716 595474
rect 345664 595410 345716 595416
rect 347780 595468 347832 595474
rect 347780 595410 347832 595416
rect 343548 588668 343600 588674
rect 343548 588610 343600 588616
rect 342904 577516 342956 577522
rect 342904 577458 342956 577464
rect 342260 516112 342312 516118
rect 342260 516054 342312 516060
rect 342272 515438 342300 516054
rect 342260 515432 342312 515438
rect 342260 515374 342312 515380
rect 342916 509182 342944 577458
rect 343560 515438 343588 588610
rect 345676 518906 345704 595410
rect 347044 588600 347096 588606
rect 347044 588542 347096 588548
rect 345848 550792 345900 550798
rect 345848 550734 345900 550740
rect 345756 549432 345808 549438
rect 345756 549374 345808 549380
rect 345664 518900 345716 518906
rect 345664 518842 345716 518848
rect 343548 515432 343600 515438
rect 343548 515374 343600 515380
rect 342904 509176 342956 509182
rect 342904 509118 342956 509124
rect 345768 506462 345796 549374
rect 345860 507686 345888 550734
rect 347056 509114 347084 588542
rect 347136 583024 347188 583030
rect 347136 582966 347188 582972
rect 347044 509108 347096 509114
rect 347044 509050 347096 509056
rect 345848 507680 345900 507686
rect 345848 507622 345900 507628
rect 347148 506462 347176 582966
rect 348424 552220 348476 552226
rect 348424 552162 348476 552168
rect 345756 506456 345808 506462
rect 345756 506398 345808 506404
rect 347136 506456 347188 506462
rect 347136 506398 347188 506404
rect 340880 505164 340932 505170
rect 340880 505106 340932 505112
rect 342168 505164 342220 505170
rect 342168 505106 342220 505112
rect 340892 505034 340920 505106
rect 340880 505028 340932 505034
rect 340880 504970 340932 504976
rect 348436 503606 348464 552162
rect 348424 503600 348476 503606
rect 348424 503542 348476 503548
rect 349816 497962 349844 641786
rect 349908 599146 349936 642194
rect 351276 639260 351328 639266
rect 351276 639202 351328 639208
rect 349896 599140 349948 599146
rect 349896 599082 349948 599088
rect 349896 589960 349948 589966
rect 349896 589902 349948 589908
rect 349908 536790 349936 589902
rect 350080 570716 350132 570722
rect 350080 570658 350132 570664
rect 349988 545760 350040 545766
rect 349988 545702 350040 545708
rect 349896 536784 349948 536790
rect 349896 536726 349948 536732
rect 349896 525088 349948 525094
rect 349896 525030 349948 525036
rect 349804 497956 349856 497962
rect 349804 497898 349856 497904
rect 349908 497593 349936 525030
rect 350000 506394 350028 545702
rect 350092 535362 350120 570658
rect 350080 535356 350132 535362
rect 350080 535298 350132 535304
rect 350540 532772 350592 532778
rect 350540 532714 350592 532720
rect 350552 532506 350580 532714
rect 350540 532500 350592 532506
rect 350540 532442 350592 532448
rect 351184 532500 351236 532506
rect 351184 532442 351236 532448
rect 350540 517608 350592 517614
rect 350540 517550 350592 517556
rect 350080 509924 350132 509930
rect 350080 509866 350132 509872
rect 349988 506388 350040 506394
rect 349988 506330 350040 506336
rect 350092 499361 350120 509866
rect 350078 499352 350134 499361
rect 350078 499287 350134 499296
rect 350092 498273 350120 499287
rect 350078 498264 350134 498273
rect 350078 498199 350134 498208
rect 349894 497584 349950 497593
rect 349894 497519 349950 497528
rect 350264 480956 350316 480962
rect 350264 480898 350316 480904
rect 338764 471980 338816 471986
rect 338764 471922 338816 471928
rect 349804 355360 349856 355366
rect 349804 355302 349856 355308
rect 346400 347812 346452 347818
rect 346400 347754 346452 347760
rect 332232 335368 332284 335374
rect 332232 335310 332284 335316
rect 327724 331560 327776 331566
rect 327724 331502 327776 331508
rect 329012 331492 329064 331498
rect 329012 331434 329064 331440
rect 327724 331356 327776 331362
rect 327724 331298 327776 331304
rect 326436 330132 326488 330138
rect 326436 330074 326488 330080
rect 326448 329868 326476 330074
rect 327736 329868 327764 331298
rect 329024 329868 329052 331434
rect 330944 331424 330996 331430
rect 330944 331366 330996 331372
rect 330956 329868 330984 331366
rect 332244 329868 332272 335310
rect 341890 332072 341946 332081
rect 341890 332007 341946 332016
rect 333520 331560 333572 331566
rect 333520 331502 333572 331508
rect 338028 331560 338080 331566
rect 338028 331502 338080 331508
rect 333532 329868 333560 331502
rect 336096 331424 336148 331430
rect 336096 331366 336148 331372
rect 334532 330064 334584 330070
rect 334532 330006 334584 330012
rect 334544 329882 334572 330006
rect 334544 329854 334834 329882
rect 336108 329868 336136 331366
rect 338040 329868 338068 331502
rect 339316 331492 339368 331498
rect 339316 331434 339368 331440
rect 339328 329868 339356 331434
rect 340236 329996 340288 330002
rect 340236 329938 340288 329944
rect 340248 329882 340276 329938
rect 340248 329854 340630 329882
rect 341904 329868 341932 332007
rect 343824 331696 343876 331702
rect 343824 331638 343876 331644
rect 343836 329868 343864 331638
rect 345112 331288 345164 331294
rect 345112 331230 345164 331236
rect 345124 329868 345152 331230
rect 346412 329868 346440 347754
rect 349712 340196 349764 340202
rect 349712 340138 349764 340144
rect 349724 332178 349752 340138
rect 349712 332172 349764 332178
rect 349712 332114 349764 332120
rect 348974 331528 349030 331537
rect 348974 331463 349030 331472
rect 347412 329928 347464 329934
rect 347464 329876 347714 329882
rect 347412 329870 347714 329876
rect 347424 329854 347714 329870
rect 348988 329868 349016 331463
rect 349816 325106 349844 355302
rect 350172 352572 350224 352578
rect 350172 352514 350224 352520
rect 349896 342916 349948 342922
rect 349896 342858 349948 342864
rect 349908 325106 349936 342858
rect 349988 332172 350040 332178
rect 349988 332114 350040 332120
rect 350000 326913 350028 332114
rect 350080 329860 350132 329866
rect 350080 329802 350132 329808
rect 349986 326904 350042 326913
rect 349986 326839 350042 326848
rect 350092 326754 350120 329802
rect 350184 327729 350212 352514
rect 350276 329089 350304 480898
rect 350356 331900 350408 331906
rect 350356 331842 350408 331848
rect 350262 329080 350318 329089
rect 350262 329015 350318 329024
rect 350170 327720 350226 327729
rect 350170 327655 350226 327664
rect 350000 326726 350120 326754
rect 350000 325694 350028 326726
rect 350000 325666 350212 325694
rect 349804 325100 349856 325106
rect 349804 325042 349856 325048
rect 349896 325100 349948 325106
rect 349896 325042 349948 325048
rect 350078 325000 350134 325009
rect 349724 324958 350078 324986
rect 347070 280634 347360 280650
rect 300124 280628 300176 280634
rect 347070 280628 347372 280634
rect 347070 280622 347320 280628
rect 300124 280570 300176 280576
rect 347320 280570 347372 280576
rect 299848 280016 299900 280022
rect 299848 279958 299900 279964
rect 300044 278254 300072 280092
rect 300032 278248 300084 278254
rect 300032 278190 300084 278196
rect 300136 223514 300164 280570
rect 301332 277982 301360 280092
rect 302252 280078 302634 280106
rect 301320 277976 301372 277982
rect 301320 277918 301372 277924
rect 301504 264240 301556 264246
rect 301504 264182 301556 264188
rect 300124 223508 300176 223514
rect 300124 223450 300176 223456
rect 299756 223100 299808 223106
rect 299756 223042 299808 223048
rect 301516 222290 301544 264182
rect 302252 223242 302280 280078
rect 303804 279948 303856 279954
rect 303804 279890 303856 279896
rect 303712 278044 303764 278050
rect 303712 277986 303764 277992
rect 302792 225820 302844 225826
rect 302792 225762 302844 225768
rect 302240 223236 302292 223242
rect 302240 223178 302292 223184
rect 301504 222284 301556 222290
rect 301504 222226 301556 222232
rect 299480 222148 299532 222154
rect 299480 222090 299532 222096
rect 300768 222148 300820 222154
rect 300768 222090 300820 222096
rect 300780 220862 300808 222090
rect 300768 220856 300820 220862
rect 300768 220798 300820 220804
rect 300780 219980 300808 220798
rect 301516 219994 301544 222226
rect 301516 219966 301806 219994
rect 302804 219980 302832 225762
rect 303724 219994 303752 277986
rect 303816 229094 303844 279890
rect 303908 278118 303936 280092
rect 305012 280078 305210 280106
rect 306668 280078 307142 280106
rect 305012 280022 305040 280078
rect 305000 280016 305052 280022
rect 305000 279958 305052 279964
rect 305644 278248 305696 278254
rect 305644 278190 305696 278196
rect 303896 278112 303948 278118
rect 303896 278054 303948 278060
rect 305000 271856 305052 271862
rect 305000 271798 305052 271804
rect 305012 229094 305040 271798
rect 303816 229066 304488 229094
rect 305012 229066 305408 229094
rect 304460 219994 304488 229066
rect 305380 219994 305408 229066
rect 305656 223582 305684 278190
rect 306668 258074 306696 280078
rect 308416 277982 308444 280092
rect 309244 280078 309718 280106
rect 310624 280078 311006 280106
rect 311912 280078 312294 280106
rect 313844 280078 314226 280106
rect 308404 277976 308456 277982
rect 308404 277918 308456 277924
rect 309140 276752 309192 276758
rect 309140 276694 309192 276700
rect 306392 258046 306696 258074
rect 305644 223576 305696 223582
rect 305644 223518 305696 223524
rect 306392 220318 306420 258046
rect 308864 227112 308916 227118
rect 308864 227054 308916 227060
rect 307852 223576 307904 223582
rect 307852 223518 307904 223524
rect 306840 223508 306892 223514
rect 306840 223450 306892 223456
rect 306380 220312 306432 220318
rect 306380 220254 306432 220260
rect 303724 219966 303830 219994
rect 304460 219966 304842 219994
rect 305380 219966 305854 219994
rect 306852 219980 306880 223450
rect 307864 219980 307892 223518
rect 308876 219980 308904 227054
rect 309152 220130 309180 276694
rect 309244 223174 309272 280078
rect 310520 279540 310572 279546
rect 310520 279482 310572 279488
rect 309232 223168 309284 223174
rect 309232 223110 309284 223116
rect 309152 220102 309456 220130
rect 309428 219994 309456 220102
rect 310532 219994 310560 279482
rect 310624 225758 310652 280078
rect 311164 275392 311216 275398
rect 311164 275334 311216 275340
rect 310612 225752 310664 225758
rect 310612 225694 310664 225700
rect 311176 223582 311204 275334
rect 311912 232558 311940 280078
rect 313280 277976 313332 277982
rect 313280 277918 313332 277924
rect 311900 232552 311952 232558
rect 311900 232494 311952 232500
rect 311164 223576 311216 223582
rect 311164 223518 311216 223524
rect 312912 223576 312964 223582
rect 312912 223518 312964 223524
rect 311900 222964 311952 222970
rect 311900 222906 311952 222912
rect 309428 219966 309902 219994
rect 310532 219966 310914 219994
rect 311912 219980 311940 222906
rect 312924 219980 312952 223518
rect 313292 220130 313320 277918
rect 313844 258074 313872 280078
rect 315500 279070 315528 280092
rect 315488 279064 315540 279070
rect 315488 279006 315540 279012
rect 316788 277982 316816 280092
rect 318076 278322 318104 280092
rect 320008 278390 320036 280092
rect 321296 279002 321324 280092
rect 321652 279472 321704 279478
rect 321652 279414 321704 279420
rect 321284 278996 321336 279002
rect 321284 278938 321336 278944
rect 319996 278384 320048 278390
rect 319996 278326 320048 278332
rect 318064 278316 318116 278322
rect 318064 278258 318116 278264
rect 317420 278044 317472 278050
rect 317420 277986 317472 277992
rect 316776 277976 316828 277982
rect 316776 277918 316828 277924
rect 314752 276752 314804 276758
rect 314752 276694 314804 276700
rect 313384 258046 313872 258074
rect 313384 221610 313412 258046
rect 314764 229094 314792 276694
rect 317432 229094 317460 277986
rect 318800 275324 318852 275330
rect 318800 275266 318852 275272
rect 318812 229094 318840 275266
rect 314764 229066 315528 229094
rect 317432 229066 317552 229094
rect 318812 229066 319576 229094
rect 314936 223236 314988 223242
rect 314936 223178 314988 223184
rect 313372 221604 313424 221610
rect 313372 221546 313424 221552
rect 313292 220102 313504 220130
rect 313476 219994 313504 220102
rect 313476 219966 313950 219994
rect 314948 219980 314976 223178
rect 315500 219994 315528 229066
rect 316960 222964 317012 222970
rect 316960 222906 317012 222912
rect 315500 219966 315974 219994
rect 316972 219980 317000 222906
rect 317524 219994 317552 229066
rect 318984 227044 319036 227050
rect 318984 226986 319036 226992
rect 317524 219966 317998 219994
rect 318996 219980 319024 226986
rect 319548 219994 319576 229066
rect 321008 223100 321060 223106
rect 321008 223042 321060 223048
rect 319548 219966 320022 219994
rect 321020 219980 321048 223042
rect 321664 219994 321692 279414
rect 322584 278458 322612 280092
rect 322572 278452 322624 278458
rect 322572 278394 322624 278400
rect 323124 277976 323176 277982
rect 323124 277918 323176 277924
rect 323136 229094 323164 277918
rect 323872 277574 323900 280092
rect 324700 280078 325174 280106
rect 323860 277568 323912 277574
rect 323860 277510 323912 277516
rect 324320 277432 324372 277438
rect 324320 277374 324372 277380
rect 324332 229094 324360 277374
rect 324700 258074 324728 280078
rect 326344 277568 326396 277574
rect 326344 277510 326396 277516
rect 324424 258046 324728 258074
rect 324424 229770 324452 258046
rect 324412 229764 324464 229770
rect 324412 229706 324464 229712
rect 325700 229764 325752 229770
rect 325700 229706 325752 229712
rect 323136 229066 323624 229094
rect 324332 229066 324728 229094
rect 323032 223168 323084 223174
rect 323032 223110 323084 223116
rect 321664 219966 322046 219994
rect 323044 219980 323072 223110
rect 323596 219994 323624 229066
rect 324700 219994 324728 229066
rect 325712 219994 325740 229706
rect 326356 223582 326384 277510
rect 327092 277438 327120 280092
rect 328012 280078 328394 280106
rect 329300 280078 329682 280106
rect 327080 277432 327132 277438
rect 327080 277374 327132 277380
rect 328012 258074 328040 280078
rect 329300 258074 329328 280078
rect 330956 278934 330984 280092
rect 332612 280078 332902 280106
rect 330944 278928 330996 278934
rect 330944 278870 330996 278876
rect 327276 258046 328040 258074
rect 328472 258046 329328 258074
rect 326344 223576 326396 223582
rect 326344 223518 326396 223524
rect 327276 219994 327304 258046
rect 328092 223100 328144 223106
rect 328092 223042 328144 223048
rect 323596 219966 324070 219994
rect 324700 219966 325082 219994
rect 325712 219966 326094 219994
rect 327106 219966 327304 219994
rect 328104 219980 328132 223042
rect 328472 220250 328500 258046
rect 332612 227118 332640 280078
rect 334176 278118 334204 280092
rect 335464 278526 335492 280092
rect 336766 280078 336964 280106
rect 335452 278520 335504 278526
rect 335452 278462 335504 278468
rect 334164 278112 334216 278118
rect 334164 278054 334216 278060
rect 335360 273964 335412 273970
rect 335360 273906 335412 273912
rect 335372 229094 335400 273906
rect 335372 229066 335768 229094
rect 332600 227112 332652 227118
rect 332600 227054 332652 227060
rect 333152 223576 333204 223582
rect 333152 223518 333204 223524
rect 329104 223168 329156 223174
rect 329104 223110 329156 223116
rect 328460 220244 328512 220250
rect 328460 220186 328512 220192
rect 329116 219980 329144 223110
rect 331128 223032 331180 223038
rect 331128 222974 331180 222980
rect 330116 222896 330168 222902
rect 330116 222838 330168 222844
rect 330128 219980 330156 222838
rect 331140 219980 331168 222974
rect 332140 222896 332192 222902
rect 332140 222838 332192 222844
rect 332152 219980 332180 222838
rect 333164 219980 333192 223518
rect 335176 223304 335228 223310
rect 335176 223246 335228 223252
rect 334164 223032 334216 223038
rect 334164 222974 334216 222980
rect 334176 219980 334204 222974
rect 335188 219980 335216 223246
rect 335740 219994 335768 229066
rect 336936 220182 336964 280078
rect 337384 278656 337436 278662
rect 337384 278598 337436 278604
rect 337200 223236 337252 223242
rect 337200 223178 337252 223184
rect 336924 220176 336976 220182
rect 336924 220118 336976 220124
rect 335740 219966 336214 219994
rect 337212 219980 337240 223178
rect 337396 221542 337424 278598
rect 338040 278458 338068 280092
rect 339972 278526 340000 280092
rect 341260 278662 341288 280092
rect 342548 278866 342576 280092
rect 342536 278860 342588 278866
rect 342536 278802 342588 278808
rect 341248 278656 341300 278662
rect 341248 278598 341300 278604
rect 339960 278520 340012 278526
rect 339960 278462 340012 278468
rect 338028 278452 338080 278458
rect 338028 278394 338080 278400
rect 338212 278112 338264 278118
rect 338212 278054 338264 278060
rect 341524 278112 341576 278118
rect 341524 278054 341576 278060
rect 337384 221536 337436 221542
rect 337384 221478 337436 221484
rect 338224 219980 338252 278054
rect 341536 223310 341564 278054
rect 343836 278050 343864 280092
rect 345768 278730 345796 280092
rect 347884 280078 348358 280106
rect 345756 278724 345808 278730
rect 345756 278666 345808 278672
rect 343824 278044 343876 278050
rect 343824 277986 343876 277992
rect 347884 260166 347912 280078
rect 349632 278798 349660 280092
rect 349620 278792 349672 278798
rect 349620 278734 349672 278740
rect 347872 260160 347924 260166
rect 347872 260102 347924 260108
rect 349724 227050 349752 324958
rect 350078 324935 350134 324944
rect 349804 324896 349856 324902
rect 349804 324838 349856 324844
rect 349896 324896 349948 324902
rect 349896 324838 349948 324844
rect 349816 315761 349844 324838
rect 349802 315752 349858 315761
rect 349802 315687 349858 315696
rect 349802 312216 349858 312225
rect 349802 312151 349858 312160
rect 349816 229770 349844 312151
rect 349908 304473 349936 324838
rect 350184 320906 350212 325666
rect 350000 320878 350212 320906
rect 350000 305833 350028 320878
rect 350368 316034 350396 331842
rect 350092 316006 350396 316034
rect 349986 305824 350042 305833
rect 349986 305759 350042 305768
rect 349894 304464 349950 304473
rect 349894 304399 349950 304408
rect 349988 303680 350040 303686
rect 349988 303622 350040 303628
rect 349804 229764 349856 229770
rect 349804 229706 349856 229712
rect 349712 227044 349764 227050
rect 349712 226986 349764 226992
rect 341524 223304 341576 223310
rect 341524 223246 341576 223252
rect 350000 223242 350028 303622
rect 350092 280634 350120 316006
rect 350080 280628 350132 280634
rect 350080 280570 350132 280576
rect 349988 223236 350040 223242
rect 349988 223178 350040 223184
rect 339224 222216 339276 222222
rect 339224 222158 339276 222164
rect 339236 219980 339264 222158
rect 341062 147520 341118 147529
rect 341062 147455 341118 147464
rect 340142 145344 340198 145353
rect 340142 145279 340198 145288
rect 340050 138680 340106 138689
rect 340050 138615 340106 138624
rect 299386 95024 299442 95033
rect 299386 94959 299442 94968
rect 299018 89040 299074 89049
rect 297364 89004 297416 89010
rect 299018 88975 299074 88984
rect 297364 88946 297416 88952
rect 296810 86048 296866 86057
rect 296810 85983 296866 85992
rect 297180 77240 297232 77246
rect 297180 77182 297232 77188
rect 297192 77081 297220 77182
rect 297178 77072 297234 77081
rect 297178 77007 297234 77016
rect 296812 73160 296864 73166
rect 296812 73102 296864 73108
rect 296824 72593 296852 73102
rect 296810 72584 296866 72593
rect 296810 72519 296866 72528
rect 297180 69012 297232 69018
rect 297180 68954 297232 68960
rect 297192 68105 297220 68954
rect 297178 68096 297234 68105
rect 297178 68031 297234 68040
rect 297376 65113 297404 88946
rect 298008 88324 298060 88330
rect 298008 88266 298060 88272
rect 298020 87553 298048 88266
rect 298006 87544 298062 87553
rect 298006 87479 298062 87488
rect 297548 85536 297600 85542
rect 297548 85478 297600 85484
rect 297560 84561 297588 85478
rect 297546 84552 297602 84561
rect 297546 84487 297602 84496
rect 297916 84176 297968 84182
rect 297916 84118 297968 84124
rect 297928 83065 297956 84118
rect 297914 83056 297970 83065
rect 297914 82991 297970 83000
rect 297916 82816 297968 82822
rect 297916 82758 297968 82764
rect 297928 81569 297956 82758
rect 297914 81560 297970 81569
rect 297914 81495 297970 81504
rect 298006 80064 298062 80073
rect 298006 79999 298008 80008
rect 298060 79999 298062 80008
rect 298008 79970 298060 79976
rect 297548 78668 297600 78674
rect 297548 78610 297600 78616
rect 297560 78577 297588 78610
rect 297546 78568 297602 78577
rect 297546 78503 297602 78512
rect 298008 75880 298060 75886
rect 298008 75822 298060 75828
rect 298020 75585 298048 75822
rect 298006 75576 298062 75585
rect 298006 75511 298062 75520
rect 298008 74520 298060 74526
rect 298008 74462 298060 74468
rect 298020 74089 298048 74462
rect 298006 74080 298062 74089
rect 298006 74015 298062 74024
rect 298008 70372 298060 70378
rect 298008 70314 298060 70320
rect 298020 69601 298048 70314
rect 298006 69592 298062 69601
rect 298006 69527 298062 69536
rect 297548 67584 297600 67590
rect 297548 67526 297600 67532
rect 297560 66609 297588 67526
rect 297546 66600 297602 66609
rect 297546 66535 297602 66544
rect 297362 65104 297418 65113
rect 297362 65039 297418 65048
rect 297916 64864 297968 64870
rect 297916 64806 297968 64812
rect 297928 63617 297956 64806
rect 297914 63608 297970 63617
rect 297914 63543 297970 63552
rect 298006 62112 298062 62121
rect 298006 62047 298008 62056
rect 298060 62047 298062 62056
rect 298008 62018 298060 62024
rect 317418 60344 317474 60353
rect 317418 60279 317474 60288
rect 296628 60240 296680 60246
rect 296628 60182 296680 60188
rect 303620 60240 303672 60246
rect 303620 60182 303672 60188
rect 303632 16574 303660 60182
rect 310520 60172 310572 60178
rect 310520 60114 310572 60120
rect 314660 60172 314712 60178
rect 314660 60114 314712 60120
rect 310532 16574 310560 60114
rect 303632 16546 303936 16574
rect 310532 16546 311480 16574
rect 296536 3800 296588 3806
rect 296536 3742 296588 3748
rect 297270 3632 297326 3641
rect 297270 3567 297326 3576
rect 300766 3632 300822 3641
rect 300766 3567 300822 3576
rect 297284 480 297312 3567
rect 300780 480 300808 3567
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 307944 3732 307996 3738
rect 307944 3674 307996 3680
rect 307956 480 307984 3674
rect 311452 480 311480 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 60114
rect 317432 16574 317460 60279
rect 340064 35358 340092 138615
rect 340156 54670 340184 145279
rect 340878 140992 340934 141001
rect 340878 140927 340934 140936
rect 340234 119232 340290 119241
rect 340234 119167 340290 119176
rect 340144 54664 340196 54670
rect 340144 54606 340196 54612
rect 340248 54534 340276 119167
rect 340326 110528 340382 110537
rect 340326 110463 340382 110472
rect 340340 57322 340368 110463
rect 340420 88732 340472 88738
rect 340420 88674 340472 88680
rect 340328 57316 340380 57322
rect 340328 57258 340380 57264
rect 340236 54528 340288 54534
rect 340236 54470 340288 54476
rect 340052 35352 340104 35358
rect 340052 35294 340104 35300
rect 317432 16546 318104 16574
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 339868 4004 339920 4010
rect 339868 3946 339920 3952
rect 332692 3936 332744 3942
rect 332692 3878 332744 3884
rect 322112 3800 322164 3806
rect 322112 3742 322164 3748
rect 325608 3800 325660 3806
rect 325608 3742 325660 3748
rect 322124 480 322152 3742
rect 325620 480 325648 3742
rect 329194 3632 329250 3641
rect 329194 3567 329250 3576
rect 329208 480 329236 3567
rect 332704 480 332732 3878
rect 336280 3868 336332 3874
rect 336280 3810 336332 3816
rect 336292 480 336320 3810
rect 339880 480 339908 3946
rect 340432 3670 340460 88674
rect 340510 75712 340566 75721
rect 340510 75647 340566 75656
rect 340524 58682 340552 75647
rect 340512 58676 340564 58682
rect 340512 58618 340564 58624
rect 340892 10334 340920 140927
rect 340970 114880 341026 114889
rect 340970 114815 341026 114824
rect 340984 18766 341012 114815
rect 341076 50386 341104 147455
rect 342258 143168 342314 143177
rect 342258 143103 342314 143112
rect 341246 132288 341302 132297
rect 341246 132223 341302 132232
rect 341154 121408 341210 121417
rect 341154 121343 341210 121352
rect 341064 50380 341116 50386
rect 341064 50322 341116 50328
rect 341168 40866 341196 121343
rect 341260 55962 341288 132223
rect 341338 112704 341394 112713
rect 341338 112639 341394 112648
rect 341352 60042 341380 112639
rect 341430 104000 341486 104009
rect 341430 103935 341486 103944
rect 341340 60036 341392 60042
rect 341340 59978 341392 59984
rect 341248 55956 341300 55962
rect 341248 55898 341300 55904
rect 341444 55894 341472 103935
rect 341522 101824 341578 101833
rect 341522 101759 341578 101768
rect 341536 57254 341564 101759
rect 341614 99648 341670 99657
rect 341614 99583 341670 99592
rect 341628 58750 341656 99583
rect 341706 97472 341762 97481
rect 341706 97407 341762 97416
rect 341720 61538 341748 97407
rect 341708 61532 341760 61538
rect 341708 61474 341760 61480
rect 341616 58744 341668 58750
rect 341616 58686 341668 58692
rect 341524 57248 341576 57254
rect 341524 57190 341576 57196
rect 341432 55888 341484 55894
rect 341432 55830 341484 55836
rect 341156 40860 341208 40866
rect 341156 40802 341208 40808
rect 340972 18760 341024 18766
rect 340972 18702 341024 18708
rect 342272 10402 342300 143103
rect 342350 136640 342406 136649
rect 342350 136575 342406 136584
rect 342364 62762 342392 136575
rect 342442 134464 342498 134473
rect 342442 134399 342498 134408
rect 342352 62756 342404 62762
rect 342352 62698 342404 62704
rect 342350 62656 342406 62665
rect 342350 62591 342406 62600
rect 342364 62150 342392 62591
rect 342352 62144 342404 62150
rect 342352 62086 342404 62092
rect 342456 57390 342484 134399
rect 342534 130112 342590 130121
rect 342534 130047 342590 130056
rect 342548 88738 342576 130047
rect 342626 127936 342682 127945
rect 342626 127871 342682 127880
rect 342536 88732 342588 88738
rect 342536 88674 342588 88680
rect 342534 80064 342590 80073
rect 342534 79999 342590 80008
rect 342444 57384 342496 57390
rect 342444 57326 342496 57332
rect 342260 10396 342312 10402
rect 342260 10338 342312 10344
rect 340880 10328 340932 10334
rect 340880 10270 340932 10276
rect 342548 4962 342576 79999
rect 342640 54602 342668 127871
rect 342718 125760 342774 125769
rect 342718 125695 342774 125704
rect 342732 61606 342760 125695
rect 342810 123584 342866 123593
rect 342810 123519 342866 123528
rect 342720 61600 342772 61606
rect 342720 61542 342772 61548
rect 342824 60110 342852 123519
rect 342904 117292 342956 117298
rect 342904 117234 342956 117240
rect 342916 117065 342944 117234
rect 342902 117056 342958 117065
rect 342902 116991 342958 117000
rect 342904 108996 342956 109002
rect 342904 108938 342956 108944
rect 342916 108361 342944 108938
rect 342902 108352 342958 108361
rect 342902 108287 342958 108296
rect 342904 106276 342956 106282
rect 342904 106218 342956 106224
rect 342916 106185 342944 106218
rect 342902 106176 342958 106185
rect 342902 106111 342958 106120
rect 343086 93120 343142 93129
rect 343086 93055 343142 93064
rect 342994 88768 343050 88777
rect 342994 88703 343050 88712
rect 342902 86592 342958 86601
rect 342902 86527 342958 86536
rect 342812 60104 342864 60110
rect 342812 60046 342864 60052
rect 342628 54596 342680 54602
rect 342628 54538 342680 54544
rect 342916 42090 342944 86527
rect 343008 61402 343036 88703
rect 343100 79393 343128 93055
rect 343178 90944 343234 90953
rect 343178 90879 343234 90888
rect 343086 79384 343142 79393
rect 343086 79319 343142 79328
rect 343086 69184 343142 69193
rect 343086 69119 343142 69128
rect 343100 69086 343128 69119
rect 343088 69080 343140 69086
rect 343088 69022 343140 69028
rect 343192 68898 343220 90879
rect 343100 68870 343220 68898
rect 343100 61470 343128 68870
rect 343178 67008 343234 67017
rect 343178 66943 343234 66952
rect 343192 66298 343220 66943
rect 343180 66292 343232 66298
rect 343180 66234 343232 66240
rect 343178 64832 343234 64841
rect 343178 64767 343234 64776
rect 343192 63578 343220 64767
rect 343180 63572 343232 63578
rect 343180 63514 343232 63520
rect 343180 62756 343232 62762
rect 343180 62698 343232 62704
rect 343088 61464 343140 61470
rect 343088 61406 343140 61412
rect 342996 61396 343048 61402
rect 342996 61338 343048 61344
rect 343192 56030 343220 62698
rect 343180 56024 343232 56030
rect 343180 55966 343232 55972
rect 346400 53100 346452 53106
rect 346400 53042 346452 53048
rect 342904 42084 342956 42090
rect 342904 42026 342956 42032
rect 346412 16574 346440 53042
rect 346412 16546 346992 16574
rect 342536 4956 342588 4962
rect 342536 4898 342588 4904
rect 340420 3664 340472 3670
rect 340420 3606 340472 3612
rect 343364 3664 343416 3670
rect 343364 3606 343416 3612
rect 343376 480 343404 3606
rect 346964 480 346992 16546
rect 350448 4956 350500 4962
rect 350448 4898 350500 4904
rect 350460 480 350488 4898
rect 350552 3942 350580 517550
rect 350816 405748 350868 405754
rect 350816 405690 350868 405696
rect 350632 400240 350684 400246
rect 350632 400182 350684 400188
rect 350644 280809 350672 400182
rect 350724 336048 350776 336054
rect 350724 335990 350776 335996
rect 350736 301889 350764 335990
rect 350722 301880 350778 301889
rect 350722 301815 350778 301824
rect 350828 299169 350856 405690
rect 350908 376780 350960 376786
rect 350908 376722 350960 376728
rect 350920 317529 350948 376722
rect 351092 334620 351144 334626
rect 351092 334562 351144 334568
rect 351000 333396 351052 333402
rect 351000 333338 351052 333344
rect 350906 317520 350962 317529
rect 350906 317455 350962 317464
rect 350906 308000 350962 308009
rect 350906 307935 350962 307944
rect 350814 299160 350870 299169
rect 350814 299095 350870 299104
rect 350722 291680 350778 291689
rect 350722 291615 350778 291624
rect 350630 280800 350686 280809
rect 350630 280735 350686 280744
rect 350736 264246 350764 291615
rect 350920 276758 350948 307935
rect 351012 284209 351040 333338
rect 351104 288289 351132 334562
rect 351090 288280 351146 288289
rect 351090 288215 351146 288224
rect 350998 284200 351054 284209
rect 350998 284135 351054 284144
rect 350908 276752 350960 276758
rect 350908 276694 350960 276700
rect 350724 264240 350776 264246
rect 350724 264182 350776 264188
rect 350540 3936 350592 3942
rect 350540 3878 350592 3884
rect 351196 3806 351224 532442
rect 351288 219434 351316 639202
rect 351380 497690 351408 642330
rect 351460 550996 351512 551002
rect 351460 550938 351512 550944
rect 351472 527134 351500 550938
rect 352472 550044 352524 550050
rect 352472 549986 352524 549992
rect 351460 527128 351512 527134
rect 351460 527070 351512 527076
rect 351460 521688 351512 521694
rect 351460 521630 351512 521636
rect 351472 498001 351500 521630
rect 352484 521626 352512 549986
rect 352472 521620 352524 521626
rect 352472 521562 352524 521568
rect 352484 521082 352512 521562
rect 352472 521076 352524 521082
rect 352472 521018 352524 521024
rect 352576 500954 352604 663750
rect 352840 662992 352892 662998
rect 352840 662934 352892 662940
rect 352656 662924 352708 662930
rect 352656 662866 352708 662872
rect 352564 500948 352616 500954
rect 352564 500890 352616 500896
rect 352564 498228 352616 498234
rect 352564 498170 352616 498176
rect 351458 497992 351514 498001
rect 351458 497927 351514 497936
rect 351368 497684 351420 497690
rect 351368 497626 351420 497632
rect 351460 429208 351512 429214
rect 351460 429150 351512 429156
rect 351368 314696 351420 314702
rect 351368 314638 351420 314644
rect 351380 222970 351408 314638
rect 351472 314129 351500 429150
rect 352104 347064 352156 347070
rect 352104 347006 352156 347012
rect 352012 334688 352064 334694
rect 352012 334630 352064 334636
rect 351918 321600 351974 321609
rect 351918 321535 351974 321544
rect 351932 314702 351960 321535
rect 351920 314696 351972 314702
rect 351920 314638 351972 314644
rect 351458 314120 351514 314129
rect 351458 314055 351514 314064
rect 351918 311400 351974 311409
rect 351918 311335 351974 311344
rect 351932 303686 351960 311335
rect 352024 306649 352052 334630
rect 352010 306640 352066 306649
rect 352010 306575 352066 306584
rect 351920 303680 351972 303686
rect 351920 303622 351972 303628
rect 351458 300520 351514 300529
rect 351458 300455 351514 300464
rect 351472 280974 351500 300455
rect 352116 297809 352144 347006
rect 352472 341556 352524 341562
rect 352472 341498 352524 341504
rect 352288 338768 352340 338774
rect 352288 338710 352340 338716
rect 352196 331492 352248 331498
rect 352196 331434 352248 331440
rect 352102 297800 352158 297809
rect 352102 297735 352158 297744
rect 351918 294400 351974 294409
rect 351918 294335 351974 294344
rect 351932 287054 351960 294335
rect 352102 293040 352158 293049
rect 352102 292975 352158 292984
rect 351932 287026 352052 287054
rect 351918 286920 351974 286929
rect 351918 286855 351974 286864
rect 351460 280968 351512 280974
rect 351460 280910 351512 280916
rect 351932 278118 351960 286855
rect 352024 281382 352052 287026
rect 352012 281376 352064 281382
rect 352012 281318 352064 281324
rect 351920 278112 351972 278118
rect 351920 278054 351972 278060
rect 352116 236706 352144 292975
rect 352208 279478 352236 331434
rect 352300 290329 352328 338710
rect 352380 333328 352432 333334
rect 352380 333270 352432 333276
rect 352392 318889 352420 333270
rect 352378 318880 352434 318889
rect 352378 318815 352434 318824
rect 352378 310040 352434 310049
rect 352378 309975 352434 309984
rect 352286 290320 352342 290329
rect 352286 290255 352342 290264
rect 352286 285560 352342 285569
rect 352286 285495 352342 285504
rect 352196 279472 352248 279478
rect 352196 279414 352248 279420
rect 352104 236700 352156 236706
rect 352104 236642 352156 236648
rect 351368 222964 351420 222970
rect 351368 222906 351420 222912
rect 352300 221474 352328 285495
rect 352392 262886 352420 309975
rect 352484 296449 352512 341498
rect 352470 296440 352526 296449
rect 352470 296375 352526 296384
rect 352380 262880 352432 262886
rect 352380 262822 352432 262828
rect 352288 221468 352340 221474
rect 352288 221410 352340 221416
rect 351276 219428 351328 219434
rect 351276 219370 351328 219376
rect 352576 60178 352604 498170
rect 352668 497622 352696 662866
rect 352748 662652 352800 662658
rect 352748 662594 352800 662600
rect 352760 497894 352788 662594
rect 352852 498166 352880 662934
rect 353024 662856 353076 662862
rect 353024 662798 353076 662804
rect 352932 662720 352984 662726
rect 352932 662662 352984 662668
rect 352840 498160 352892 498166
rect 352840 498102 352892 498108
rect 352748 497888 352800 497894
rect 352748 497830 352800 497836
rect 352944 497826 352972 662662
rect 353036 520266 353064 662798
rect 355324 662788 355376 662794
rect 355324 662730 355376 662736
rect 353116 656940 353168 656946
rect 353116 656882 353168 656888
rect 353128 599078 353156 656882
rect 353208 642728 353260 642734
rect 353208 642670 353260 642676
rect 353220 599214 353248 642670
rect 354036 639328 354088 639334
rect 354036 639270 354088 639276
rect 353944 639192 353996 639198
rect 353944 639134 353996 639140
rect 353208 599208 353260 599214
rect 353208 599150 353260 599156
rect 353116 599072 353168 599078
rect 353116 599014 353168 599020
rect 353116 584452 353168 584458
rect 353116 584394 353168 584400
rect 353128 535294 353156 584394
rect 353208 549500 353260 549506
rect 353208 549442 353260 549448
rect 353116 535288 353168 535294
rect 353116 535230 353168 535236
rect 353116 520328 353168 520334
rect 353116 520270 353168 520276
rect 353024 520260 353076 520266
rect 353024 520202 353076 520208
rect 353024 515432 353076 515438
rect 353024 515374 353076 515380
rect 353036 499322 353064 515374
rect 353128 500886 353156 520270
rect 353220 509250 353248 549442
rect 353482 530632 353538 530641
rect 353482 530567 353538 530576
rect 353300 521076 353352 521082
rect 353300 521018 353352 521024
rect 353208 509244 353260 509250
rect 353208 509186 353260 509192
rect 353116 500880 353168 500886
rect 353116 500822 353168 500828
rect 353024 499316 353076 499322
rect 353024 499258 353076 499264
rect 353036 498234 353064 499258
rect 353024 498228 353076 498234
rect 353024 498170 353076 498176
rect 352932 497820 352984 497826
rect 352932 497762 352984 497768
rect 352656 497616 352708 497622
rect 352656 497558 352708 497564
rect 352656 354000 352708 354006
rect 352656 353942 352708 353948
rect 352668 282849 352696 353942
rect 352746 323640 352802 323649
rect 352746 323575 352802 323584
rect 352654 282840 352710 282849
rect 352654 282775 352710 282784
rect 352760 261526 352788 323575
rect 352748 261520 352800 261526
rect 352748 261462 352800 261468
rect 352564 60172 352616 60178
rect 352564 60114 352616 60120
rect 351184 3800 351236 3806
rect 351184 3742 351236 3748
rect 353312 3670 353340 521018
rect 353392 498908 353444 498914
rect 353392 498850 353444 498856
rect 353404 4010 353432 498850
rect 353496 291689 353524 530567
rect 353576 331560 353628 331566
rect 353576 331502 353628 331508
rect 353482 291680 353538 291689
rect 353482 291615 353538 291624
rect 353588 223106 353616 331502
rect 353668 331356 353720 331362
rect 353668 331298 353720 331304
rect 353576 223100 353628 223106
rect 353576 223042 353628 223048
rect 353680 222902 353708 331298
rect 353668 222896 353720 222902
rect 353668 222838 353720 222844
rect 353956 139398 353984 639134
rect 354048 313274 354076 639270
rect 355232 557048 355284 557054
rect 355232 556990 355284 556996
rect 354956 552288 355008 552294
rect 354956 552230 355008 552236
rect 354220 551132 354272 551138
rect 354220 551074 354272 551080
rect 354128 541680 354180 541686
rect 354128 541622 354180 541628
rect 354140 497350 354168 541622
rect 354232 529922 354260 551074
rect 354968 543734 354996 552230
rect 355140 550112 355192 550118
rect 355140 550054 355192 550060
rect 355048 549976 355100 549982
rect 355048 549918 355100 549924
rect 355060 546802 355088 549918
rect 355152 549370 355180 550054
rect 355140 549364 355192 549370
rect 355140 549306 355192 549312
rect 355060 546774 355180 546802
rect 354968 543706 355088 543734
rect 354220 529916 354272 529922
rect 354220 529858 354272 529864
rect 355060 525774 355088 543706
rect 355152 532710 355180 546774
rect 355140 532704 355192 532710
rect 355140 532646 355192 532652
rect 355244 532506 355272 556990
rect 355232 532500 355284 532506
rect 355232 532442 355284 532448
rect 355336 527134 355364 662730
rect 355428 536722 355456 663818
rect 356888 661496 356940 661502
rect 356888 661438 356940 661444
rect 355968 642388 356020 642394
rect 355968 642330 356020 642336
rect 355600 642184 355652 642190
rect 355600 642126 355652 642132
rect 355508 640960 355560 640966
rect 355508 640902 355560 640908
rect 355520 598806 355548 640902
rect 355612 599282 355640 642126
rect 355600 599276 355652 599282
rect 355600 599218 355652 599224
rect 355508 598800 355560 598806
rect 355508 598742 355560 598748
rect 355876 567860 355928 567866
rect 355876 567802 355928 567808
rect 355888 557534 355916 567802
rect 355612 557506 355916 557534
rect 355508 550928 355560 550934
rect 355508 550870 355560 550876
rect 355416 536716 355468 536722
rect 355416 536658 355468 536664
rect 355324 527128 355376 527134
rect 355324 527070 355376 527076
rect 355048 525768 355100 525774
rect 355048 525710 355100 525716
rect 355416 519580 355468 519586
rect 355416 519522 355468 519528
rect 355324 513392 355376 513398
rect 355324 513334 355376 513340
rect 355336 499574 355364 513334
rect 355244 499546 355364 499574
rect 355244 498953 355272 499546
rect 355230 498944 355286 498953
rect 355230 498879 355286 498888
rect 354128 497344 354180 497350
rect 354128 497286 354180 497292
rect 355244 489914 355272 498879
rect 355428 498166 355456 519522
rect 355520 507822 355548 550870
rect 355612 550866 355640 557506
rect 355692 554124 355744 554130
rect 355692 554066 355744 554072
rect 355600 550860 355652 550866
rect 355600 550802 355652 550808
rect 355612 510610 355640 550802
rect 355704 513330 355732 554066
rect 355784 552356 355836 552362
rect 355784 552298 355836 552304
rect 355796 522986 355824 552298
rect 355876 523048 355928 523054
rect 355876 522990 355928 522996
rect 355784 522980 355836 522986
rect 355784 522922 355836 522928
rect 355692 513324 355744 513330
rect 355692 513266 355744 513272
rect 355600 510604 355652 510610
rect 355600 510546 355652 510552
rect 355508 507816 355560 507822
rect 355508 507758 355560 507764
rect 355508 502376 355560 502382
rect 355508 502318 355560 502324
rect 355324 498160 355376 498166
rect 355324 498102 355376 498108
rect 355416 498160 355468 498166
rect 355416 498102 355468 498108
rect 355336 497758 355364 498102
rect 355324 497752 355376 497758
rect 355324 497694 355376 497700
rect 355244 489886 355364 489914
rect 354680 331424 354732 331430
rect 354680 331366 354732 331372
rect 354036 313268 354088 313274
rect 354036 313210 354088 313216
rect 354692 223174 354720 331366
rect 354772 331288 354824 331294
rect 354772 331230 354824 331236
rect 354680 223168 354732 223174
rect 354680 223110 354732 223116
rect 354784 223038 354812 331230
rect 354772 223032 354824 223038
rect 354772 222974 354824 222980
rect 353944 139392 353996 139398
rect 353944 139334 353996 139340
rect 353576 13116 353628 13122
rect 353576 13058 353628 13064
rect 353392 4004 353444 4010
rect 353392 3946 353444 3952
rect 353300 3664 353352 3670
rect 353300 3606 353352 3612
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 13058
rect 355336 3738 355364 489886
rect 355428 3874 355456 498102
rect 355520 497865 355548 502318
rect 355506 497856 355562 497865
rect 355506 497791 355562 497800
rect 355888 497457 355916 522990
rect 355980 499526 356008 642330
rect 356796 640620 356848 640626
rect 356796 640562 356848 640568
rect 356704 640552 356756 640558
rect 356704 640494 356756 640500
rect 356060 552424 356112 552430
rect 356060 552366 356112 552372
rect 356072 548622 356100 552366
rect 356060 548616 356112 548622
rect 356060 548558 356112 548564
rect 356612 505776 356664 505782
rect 356612 505718 356664 505724
rect 355968 499520 356020 499526
rect 355968 499462 356020 499468
rect 356624 498982 356652 505718
rect 356612 498976 356664 498982
rect 356612 498918 356664 498924
rect 355874 497448 355930 497457
rect 355874 497383 355930 497392
rect 356716 60722 356744 640494
rect 356808 259418 356836 640562
rect 356900 553042 356928 661438
rect 356980 659932 357032 659938
rect 356980 659874 357032 659880
rect 356888 553036 356940 553042
rect 356888 552978 356940 552984
rect 356992 552974 357020 659874
rect 357348 642864 357400 642870
rect 357348 642806 357400 642812
rect 357256 642660 357308 642666
rect 357256 642602 357308 642608
rect 357072 641912 357124 641918
rect 357072 641854 357124 641860
rect 357084 599418 357112 641854
rect 357164 640892 357216 640898
rect 357164 640834 357216 640840
rect 357072 599412 357124 599418
rect 357072 599354 357124 599360
rect 357176 598670 357204 640834
rect 357164 598664 357216 598670
rect 357164 598606 357216 598612
rect 357072 598528 357124 598534
rect 357072 598470 357124 598476
rect 356980 552968 357032 552974
rect 356980 552910 357032 552916
rect 356980 550656 357032 550662
rect 356980 550598 357032 550604
rect 356888 550180 356940 550186
rect 356888 550122 356940 550128
rect 356900 517614 356928 550122
rect 356992 528562 357020 550598
rect 356980 528556 357032 528562
rect 356980 528498 357032 528504
rect 356888 517608 356940 517614
rect 356888 517550 356940 517556
rect 356888 516724 356940 516730
rect 356888 516666 356940 516672
rect 356900 497321 356928 516666
rect 356980 511284 357032 511290
rect 356980 511226 357032 511232
rect 356992 498778 357020 511226
rect 357084 499050 357112 598470
rect 357164 573368 357216 573374
rect 357164 573310 357216 573316
rect 357176 550361 357204 573310
rect 357162 550352 357218 550361
rect 357162 550287 357218 550296
rect 357162 516216 357218 516225
rect 357162 516151 357218 516160
rect 357176 512650 357204 516151
rect 357164 512644 357216 512650
rect 357164 512586 357216 512592
rect 357164 507884 357216 507890
rect 357164 507826 357216 507832
rect 357176 499497 357204 507826
rect 357162 499488 357218 499497
rect 357162 499423 357218 499432
rect 357072 499044 357124 499050
rect 357072 498986 357124 498992
rect 356980 498772 357032 498778
rect 356980 498714 357032 498720
rect 357268 498030 357296 642602
rect 357360 498098 357388 642806
rect 359464 642592 359516 642598
rect 359464 642534 359516 642540
rect 358820 641776 358872 641782
rect 358820 641718 358872 641724
rect 358544 641232 358596 641238
rect 358544 641174 358596 641180
rect 357808 640824 357860 640830
rect 357808 640766 357860 640772
rect 357622 548584 357678 548593
rect 357622 548519 357678 548528
rect 357440 547868 357492 547874
rect 357440 547810 357492 547816
rect 357452 547777 357480 547810
rect 357438 547768 357494 547777
rect 357438 547703 357494 547712
rect 357440 546440 357492 546446
rect 357440 546382 357492 546388
rect 357452 546009 357480 546382
rect 357438 546000 357494 546009
rect 357438 545935 357494 545944
rect 357440 545080 357492 545086
rect 357440 545022 357492 545028
rect 357452 544649 357480 545022
rect 357438 544640 357494 544649
rect 357438 544575 357494 544584
rect 357530 543552 357586 543561
rect 357530 543487 357586 543496
rect 357544 543046 357572 543487
rect 357532 543040 357584 543046
rect 357532 542982 357584 542988
rect 357440 539572 357492 539578
rect 357440 539514 357492 539520
rect 357452 539209 357480 539514
rect 357438 539200 357494 539209
rect 357438 539135 357494 539144
rect 357440 536784 357492 536790
rect 357438 536752 357440 536761
rect 357492 536752 357494 536761
rect 357438 536687 357494 536696
rect 357440 535424 357492 535430
rect 357438 535392 357440 535401
rect 357492 535392 357494 535401
rect 357438 535327 357494 535336
rect 357532 535356 357584 535362
rect 357532 535298 357584 535304
rect 357440 535288 357492 535294
rect 357440 535230 357492 535236
rect 357452 534993 357480 535230
rect 357438 534984 357494 534993
rect 357438 534919 357494 534928
rect 357544 534585 357572 535298
rect 357530 534576 357586 534585
rect 357530 534511 357586 534520
rect 357440 532636 357492 532642
rect 357440 532578 357492 532584
rect 357452 532409 357480 532578
rect 357532 532568 357584 532574
rect 357532 532510 357584 532516
rect 357438 532400 357494 532409
rect 357438 532335 357494 532344
rect 357544 531865 357572 532510
rect 357530 531856 357586 531865
rect 357530 531791 357586 531800
rect 357440 529848 357492 529854
rect 357440 529790 357492 529796
rect 357452 529553 357480 529790
rect 357438 529544 357494 529553
rect 357438 529479 357494 529488
rect 357440 527060 357492 527066
rect 357440 527002 357492 527008
rect 357452 526833 357480 527002
rect 357438 526824 357494 526833
rect 357438 526759 357494 526768
rect 357440 524408 357492 524414
rect 357440 524350 357492 524356
rect 357452 523705 357480 524350
rect 357438 523696 357494 523705
rect 357438 523631 357494 523640
rect 357636 522986 357664 548519
rect 357716 533384 357768 533390
rect 357714 533352 357716 533361
rect 357768 533352 357770 533361
rect 357714 533287 357770 533296
rect 357716 530324 357768 530330
rect 357716 530266 357768 530272
rect 357624 522980 357676 522986
rect 357624 522922 357676 522928
rect 357440 520260 357492 520266
rect 357440 520202 357492 520208
rect 357452 519625 357480 520202
rect 357438 519616 357494 519625
rect 357438 519551 357494 519560
rect 357440 518900 357492 518906
rect 357440 518842 357492 518848
rect 357452 518809 357480 518842
rect 357438 518800 357494 518809
rect 357438 518735 357494 518744
rect 357530 517576 357586 517585
rect 357530 517511 357532 517520
rect 357584 517511 357586 517520
rect 357532 517482 357584 517488
rect 357440 517472 357492 517478
rect 357438 517440 357440 517449
rect 357492 517440 357494 517449
rect 357438 517375 357494 517384
rect 357440 514752 357492 514758
rect 357438 514720 357440 514729
rect 357492 514720 357494 514729
rect 357438 514655 357494 514664
rect 357440 513256 357492 513262
rect 357440 513198 357492 513204
rect 357452 512825 357480 513198
rect 357438 512816 357494 512825
rect 357438 512751 357494 512760
rect 357440 511964 357492 511970
rect 357440 511906 357492 511912
rect 357452 511465 357480 511906
rect 357622 511592 357678 511601
rect 357622 511527 357678 511536
rect 357438 511456 357494 511465
rect 357438 511391 357494 511400
rect 357440 510536 357492 510542
rect 357440 510478 357492 510484
rect 357452 510377 357480 510478
rect 357438 510368 357494 510377
rect 357438 510303 357494 510312
rect 357532 509176 357584 509182
rect 357532 509118 357584 509124
rect 357440 509108 357492 509114
rect 357440 509050 357492 509056
rect 357452 509017 357480 509050
rect 357438 509008 357494 509017
rect 357438 508943 357494 508952
rect 357544 508745 357572 509118
rect 357530 508736 357586 508745
rect 357530 508671 357586 508680
rect 357440 507748 357492 507754
rect 357440 507690 357492 507696
rect 357452 507385 357480 507690
rect 357438 507376 357494 507385
rect 357438 507311 357494 507320
rect 357440 506456 357492 506462
rect 357440 506398 357492 506404
rect 357452 506297 357480 506398
rect 357532 506388 357584 506394
rect 357532 506330 357584 506336
rect 357438 506288 357494 506297
rect 357438 506223 357494 506232
rect 357544 505889 357572 506330
rect 357530 505880 357586 505889
rect 357530 505815 357586 505824
rect 357440 505096 357492 505102
rect 357440 505038 357492 505044
rect 357452 504665 357480 505038
rect 357438 504656 357494 504665
rect 357438 504591 357494 504600
rect 357440 503668 357492 503674
rect 357440 503610 357492 503616
rect 357452 503305 357480 503610
rect 357438 503296 357494 503305
rect 357438 503231 357494 503240
rect 357440 502308 357492 502314
rect 357440 502250 357492 502256
rect 357452 501945 357480 502250
rect 357438 501936 357494 501945
rect 357438 501871 357494 501880
rect 357348 498092 357400 498098
rect 357348 498034 357400 498040
rect 357256 498024 357308 498030
rect 357256 497966 357308 497972
rect 356886 497312 356942 497321
rect 356886 497247 356942 497256
rect 356796 259412 356848 259418
rect 356796 259354 356848 259360
rect 356704 60716 356756 60722
rect 356704 60658 356756 60664
rect 357440 17264 357492 17270
rect 357440 17206 357492 17212
rect 357452 16574 357480 17206
rect 357452 16546 357572 16574
rect 355416 3868 355468 3874
rect 355416 3810 355468 3816
rect 355324 3732 355376 3738
rect 355324 3674 355376 3680
rect 357544 480 357572 16546
rect 357636 5030 357664 511527
rect 357728 509234 357756 530266
rect 357820 510105 357848 640766
rect 357900 640552 357952 640558
rect 357900 640494 357952 640500
rect 357912 548457 357940 640494
rect 358452 639668 358504 639674
rect 358452 639610 358504 639616
rect 358176 566568 358228 566574
rect 358176 566510 358228 566516
rect 358084 562488 358136 562494
rect 358084 562430 358136 562436
rect 357898 548448 357954 548457
rect 357898 548383 357954 548392
rect 358096 543734 358124 562430
rect 358004 543706 358124 543734
rect 358004 543561 358032 543706
rect 357990 543552 358046 543561
rect 357990 543487 358046 543496
rect 357900 536716 357952 536722
rect 357900 536658 357952 536664
rect 357912 536625 357940 536658
rect 357898 536616 357954 536625
rect 357898 536551 357954 536560
rect 358188 533526 358216 566510
rect 358268 559632 358320 559638
rect 358268 559574 358320 559580
rect 358176 533520 358228 533526
rect 358176 533462 358228 533468
rect 358280 533406 358308 559574
rect 358360 556844 358412 556850
rect 358360 556786 358412 556792
rect 358372 538121 358400 556786
rect 358464 540977 358492 639610
rect 358450 540968 358506 540977
rect 358450 540903 358506 540912
rect 358358 538112 358414 538121
rect 358358 538047 358414 538056
rect 358372 536858 358400 538047
rect 358360 536852 358412 536858
rect 358360 536794 358412 536800
rect 358004 533378 358308 533406
rect 357900 527128 357952 527134
rect 357900 527070 357952 527076
rect 357912 526425 357940 527070
rect 357898 526416 357954 526425
rect 357898 526351 357954 526360
rect 358004 521937 358032 533378
rect 358174 528592 358230 528601
rect 358174 528527 358230 528536
rect 358082 525192 358138 525201
rect 358082 525127 358138 525136
rect 357990 521928 358046 521937
rect 357990 521863 358046 521872
rect 358096 514894 358124 525127
rect 358084 514888 358136 514894
rect 358084 514830 358136 514836
rect 357806 510096 357862 510105
rect 357806 510031 357862 510040
rect 357728 509206 357848 509234
rect 357820 507793 357848 509206
rect 357806 507784 357862 507793
rect 357806 507719 357862 507728
rect 358188 496806 358216 528527
rect 358266 519752 358322 519761
rect 358266 519687 358322 519696
rect 358280 513330 358308 519687
rect 358268 513324 358320 513330
rect 358268 513266 358320 513272
rect 358266 513224 358322 513233
rect 358266 513159 358322 513168
rect 358176 496800 358228 496806
rect 358176 496742 358228 496748
rect 358280 494018 358308 513159
rect 358372 500818 358400 536794
rect 358556 527785 358584 641174
rect 358636 639600 358688 639606
rect 358636 639542 358688 639548
rect 358542 527776 358598 527785
rect 358542 527711 358598 527720
rect 358542 526960 358598 526969
rect 358542 526895 358598 526904
rect 358450 522064 358506 522073
rect 358450 521999 358506 522008
rect 358360 500812 358412 500818
rect 358360 500754 358412 500760
rect 358268 494012 358320 494018
rect 358268 493954 358320 493960
rect 358464 177342 358492 521999
rect 358556 516225 358584 526895
rect 358648 525065 358676 639542
rect 358728 553444 358780 553450
rect 358728 553386 358780 553392
rect 358740 545057 358768 553386
rect 358726 545048 358782 545057
rect 358726 544983 358782 544992
rect 358832 543425 358860 641718
rect 359188 640756 359240 640762
rect 359188 640698 359240 640704
rect 358912 639396 358964 639402
rect 358912 639338 358964 639344
rect 358818 543416 358874 543425
rect 358818 543351 358874 543360
rect 358818 539336 358874 539345
rect 358818 539271 358874 539280
rect 358634 525056 358690 525065
rect 358634 524991 358690 525000
rect 358634 523832 358690 523841
rect 358634 523767 358690 523776
rect 358542 516216 358598 516225
rect 358542 516151 358598 516160
rect 358542 515128 358598 515137
rect 358542 515063 358598 515072
rect 358452 177336 358504 177342
rect 358452 177278 358504 177284
rect 358556 89078 358584 515063
rect 358544 89072 358596 89078
rect 358544 89014 358596 89020
rect 358648 89010 358676 523767
rect 358728 507884 358780 507890
rect 358728 507826 358780 507832
rect 358740 503713 358768 507826
rect 358726 503704 358782 503713
rect 358726 503639 358782 503648
rect 358636 89004 358688 89010
rect 358636 88946 358688 88952
rect 358832 86970 358860 539271
rect 358924 537849 358952 639338
rect 359096 563712 359148 563718
rect 359096 563654 359148 563660
rect 359004 558340 359056 558346
rect 359004 558282 359056 558288
rect 358910 537840 358966 537849
rect 358910 537775 358966 537784
rect 358910 532808 358966 532817
rect 358910 532743 358966 532752
rect 358924 489190 358952 532743
rect 359016 513369 359044 558282
rect 359108 521665 359136 563654
rect 359200 542337 359228 640698
rect 359372 556912 359424 556918
rect 359372 556854 359424 556860
rect 359280 555552 359332 555558
rect 359280 555494 359332 555500
rect 359186 542328 359242 542337
rect 359186 542263 359242 542272
rect 359094 521656 359150 521665
rect 359094 521591 359150 521600
rect 359292 520985 359320 555494
rect 359384 528329 359412 556854
rect 359476 530330 359504 642534
rect 359740 641980 359792 641986
rect 359740 641922 359792 641928
rect 359648 599208 359700 599214
rect 359648 599150 359700 599156
rect 359660 598942 359688 599150
rect 359648 598936 359700 598942
rect 359648 598878 359700 598884
rect 359752 538214 359780 641922
rect 360108 641844 360160 641850
rect 360108 641786 360160 641792
rect 360016 640484 360068 640490
rect 360016 640426 360068 640432
rect 360028 599214 360056 640426
rect 360016 599208 360068 599214
rect 360016 599150 360068 599156
rect 360120 553110 360148 641786
rect 360108 553104 360160 553110
rect 360108 553046 360160 553052
rect 360660 552832 360712 552838
rect 360660 552774 360712 552780
rect 360108 551540 360160 551546
rect 360108 551482 360160 551488
rect 360120 549930 360148 551482
rect 360042 549902 360148 549930
rect 360672 549916 360700 552774
rect 360856 550633 360884 700402
rect 397472 698970 397500 703520
rect 406384 700324 406436 700330
rect 406384 700266 406436 700272
rect 397460 698964 397512 698970
rect 397460 698906 397512 698912
rect 403716 670744 403768 670750
rect 403716 670686 403768 670692
rect 401600 661428 401652 661434
rect 401600 661370 401652 661376
rect 401612 661337 401640 661370
rect 401598 661328 401654 661337
rect 401598 661263 401654 661272
rect 371700 642864 371752 642870
rect 371700 642806 371752 642812
rect 361028 642796 361080 642802
rect 361028 642738 361080 642744
rect 360934 641880 360990 641889
rect 360934 641815 360990 641824
rect 360948 551993 360976 641815
rect 361040 599010 361068 642738
rect 370044 642524 370096 642530
rect 370044 642466 370096 642472
rect 361764 642456 361816 642462
rect 361764 642398 361816 642404
rect 366180 642456 366232 642462
rect 366180 642398 366232 642404
rect 361212 640416 361264 640422
rect 361212 640358 361264 640364
rect 361120 640348 361172 640354
rect 361120 640290 361172 640296
rect 361028 599004 361080 599010
rect 361028 598946 361080 598952
rect 361132 598738 361160 640290
rect 361224 598874 361252 640358
rect 361776 639962 361804 642398
rect 365536 642320 365588 642326
rect 365074 642288 365130 642297
rect 365536 642262 365588 642268
rect 365074 642223 365130 642232
rect 363420 642048 363472 642054
rect 363420 641990 363472 641996
rect 361946 639976 362002 639985
rect 361776 639948 361946 639962
rect 361790 639934 361946 639948
rect 363432 639948 363460 641990
rect 364550 639946 364840 639962
rect 365088 639948 365116 642223
rect 365548 640121 365576 642262
rect 365534 640112 365590 640121
rect 365534 640047 365590 640056
rect 366192 639948 366220 642398
rect 368938 642016 368994 642025
rect 368938 641951 368994 641960
rect 368388 641844 368440 641850
rect 368388 641786 368440 641792
rect 366732 641776 366784 641782
rect 366732 641718 366784 641724
rect 366744 639948 366772 641718
rect 367560 640008 367612 640014
rect 367310 639956 367560 639962
rect 367310 639950 367612 639956
rect 364550 639940 364852 639946
rect 364550 639934 364800 639940
rect 361946 639911 362002 639920
rect 367310 639934 367600 639950
rect 368400 639948 368428 641786
rect 368952 639948 368980 641951
rect 369490 641744 369546 641753
rect 369490 641679 369546 641688
rect 369504 639948 369532 641679
rect 370056 639948 370084 642466
rect 371148 642116 371200 642122
rect 371148 642058 371200 642064
rect 371160 639948 371188 642058
rect 371712 639948 371740 642806
rect 379980 642796 380032 642802
rect 379980 642738 380032 642744
rect 376116 642592 376168 642598
rect 376116 642534 376168 642540
rect 376208 642592 376260 642598
rect 376208 642534 376260 642540
rect 374460 642048 374512 642054
rect 374460 641990 374512 641996
rect 373356 641980 373408 641986
rect 373356 641922 373408 641928
rect 373368 639948 373396 641922
rect 374472 639948 374500 641990
rect 375564 641776 375616 641782
rect 375564 641718 375616 641724
rect 375576 639948 375604 641718
rect 376128 639948 376156 642534
rect 376220 641782 376248 642534
rect 377772 642252 377824 642258
rect 377772 642194 377824 642200
rect 376208 641776 376260 641782
rect 376208 641718 376260 641724
rect 377784 639948 377812 642194
rect 378048 641844 378100 641850
rect 378048 641786 378100 641792
rect 378060 640937 378088 641786
rect 378324 640960 378376 640966
rect 378046 640928 378102 640937
rect 378324 640902 378376 640908
rect 378046 640863 378102 640872
rect 378336 639948 378364 640902
rect 379428 640484 379480 640490
rect 379428 640426 379480 640432
rect 379440 639948 379468 640426
rect 379992 639948 380020 642738
rect 382188 642728 382240 642734
rect 382188 642670 382240 642676
rect 381084 641912 381136 641918
rect 381084 641854 381136 641860
rect 381096 639948 381124 641854
rect 382200 639948 382228 642670
rect 388812 642660 388864 642666
rect 388812 642602 388864 642608
rect 392676 642660 392728 642666
rect 392676 642602 392728 642608
rect 399300 642660 399352 642666
rect 399300 642602 399352 642608
rect 383292 642320 383344 642326
rect 383292 642262 383344 642268
rect 383304 639948 383332 642262
rect 387156 642252 387208 642258
rect 387156 642194 387208 642200
rect 386052 642184 386104 642190
rect 386052 642126 386104 642132
rect 383844 640892 383896 640898
rect 383844 640834 383896 640840
rect 383856 639948 383884 640834
rect 384948 640688 385000 640694
rect 384948 640630 385000 640636
rect 384396 640416 384448 640422
rect 384396 640358 384448 640364
rect 384408 639948 384436 640358
rect 384960 639948 384988 640630
rect 385500 640348 385552 640354
rect 385500 640290 385552 640296
rect 385512 639948 385540 640290
rect 386064 639948 386092 642126
rect 386604 641844 386656 641850
rect 386604 641786 386656 641792
rect 386616 639948 386644 641786
rect 387168 639948 387196 642194
rect 388260 640824 388312 640830
rect 388260 640766 388312 640772
rect 387708 640688 387760 640694
rect 387708 640630 387760 640636
rect 387720 639948 387748 640630
rect 388272 639948 388300 640766
rect 388824 639948 388852 642602
rect 391020 642388 391072 642394
rect 391020 642330 391072 642336
rect 392124 642388 392176 642394
rect 392124 642330 392176 642336
rect 390466 642152 390522 642161
rect 390466 642087 390522 642096
rect 389364 640756 389416 640762
rect 389364 640698 389416 640704
rect 389376 639948 389404 640698
rect 389916 640620 389968 640626
rect 389916 640562 389968 640568
rect 389928 639948 389956 640562
rect 390480 639948 390508 642087
rect 391032 639948 391060 642330
rect 391572 641232 391624 641238
rect 391572 641174 391624 641180
rect 391584 639948 391612 641174
rect 392136 639948 392164 642330
rect 392688 639948 392716 642602
rect 399116 642456 399168 642462
rect 399116 642398 399168 642404
rect 393228 642320 393280 642326
rect 393228 642262 393280 642268
rect 393240 639948 393268 642262
rect 394332 642184 394384 642190
rect 394332 642126 394384 642132
rect 393780 641844 393832 641850
rect 393780 641786 393832 641792
rect 393792 639948 393820 641786
rect 394344 639948 394372 642126
rect 394884 641912 394936 641918
rect 394884 641854 394936 641860
rect 397090 641880 397146 641889
rect 394896 639948 394924 641854
rect 397090 641815 397146 641824
rect 395436 641776 395488 641782
rect 395436 641718 395488 641724
rect 395448 639948 395476 641718
rect 396540 640552 396592 640558
rect 396540 640494 396592 640500
rect 396552 639948 396580 640494
rect 397104 639948 397132 641815
rect 398470 641744 398526 641753
rect 398470 641679 398526 641688
rect 398484 641170 398512 641679
rect 398472 641164 398524 641170
rect 398472 641106 398524 641112
rect 398484 639962 398512 641106
rect 373264 639940 373316 639946
rect 364800 639882 364852 639888
rect 398222 639934 398972 639962
rect 373264 639882 373316 639888
rect 365720 639872 365772 639878
rect 365654 639820 365720 639826
rect 373172 639872 373224 639878
rect 365654 639814 365772 639820
rect 365654 639798 365760 639814
rect 367862 639810 368152 639826
rect 373172 639814 373224 639820
rect 367862 639804 368164 639810
rect 367862 639798 368112 639804
rect 368112 639746 368164 639752
rect 372344 639804 372396 639810
rect 372344 639746 372396 639752
rect 362590 639568 362646 639577
rect 362646 639526 362894 639554
rect 362590 639503 362646 639512
rect 362590 639432 362646 639441
rect 362342 639390 362590 639418
rect 364062 639432 364118 639441
rect 363998 639390 364062 639418
rect 362590 639367 362646 639376
rect 371896 639402 372278 639418
rect 372356 639402 372384 639746
rect 372830 639402 373120 639418
rect 373184 639402 373212 639814
rect 373276 639402 373304 639882
rect 382372 639736 382424 639742
rect 374656 639674 375038 639690
rect 374644 639668 375038 639674
rect 374696 639662 375038 639668
rect 377246 639674 377536 639690
rect 382424 639684 382766 639690
rect 382372 639678 382766 639684
rect 377246 639668 377548 639674
rect 377246 639662 377496 639668
rect 374644 639610 374696 639616
rect 382384 639662 382766 639678
rect 377496 639610 377548 639616
rect 376300 639600 376352 639606
rect 385684 639600 385736 639606
rect 381266 639568 381322 639577
rect 376352 639548 376694 639554
rect 376300 639542 376694 639548
rect 376312 639526 376694 639542
rect 378520 639538 378902 639554
rect 378508 639532 378902 639538
rect 378560 639526 378902 639532
rect 385736 639560 385908 639588
rect 385684 639542 385736 639548
rect 385880 639554 385908 639560
rect 386142 639568 386198 639577
rect 385880 639526 386000 639554
rect 381266 639503 381322 639512
rect 378508 639474 378560 639480
rect 380164 639464 380216 639470
rect 373934 639402 374040 639418
rect 380216 639412 380558 639418
rect 380164 639406 380558 639412
rect 364062 639367 364118 639376
rect 371884 639396 372278 639402
rect 371936 639390 372278 639396
rect 372344 639396 372396 639402
rect 371884 639338 371936 639344
rect 372830 639396 373132 639402
rect 372830 639390 373080 639396
rect 372344 639338 372396 639344
rect 373080 639338 373132 639344
rect 373172 639396 373224 639402
rect 373172 639338 373224 639344
rect 373264 639396 373316 639402
rect 373934 639396 374052 639402
rect 373934 639390 374000 639396
rect 373264 639338 373316 639344
rect 380176 639390 380558 639406
rect 381280 639402 381308 639503
rect 381358 639432 381414 639441
rect 381268 639396 381320 639402
rect 374000 639338 374052 639344
rect 381726 639432 381782 639441
rect 381414 639390 381662 639418
rect 381358 639367 381414 639376
rect 381726 639367 381728 639376
rect 381268 639338 381320 639344
rect 381780 639367 381782 639376
rect 385866 639432 385922 639441
rect 385972 639402 386000 639526
rect 386142 639503 386198 639512
rect 386156 639402 386184 639503
rect 396264 639464 396316 639470
rect 396014 639412 396264 639418
rect 396014 639406 396316 639412
rect 385866 639367 385868 639376
rect 381728 639338 381780 639344
rect 385920 639367 385922 639376
rect 385960 639396 386012 639402
rect 385868 639338 385920 639344
rect 385960 639338 386012 639344
rect 386144 639396 386196 639402
rect 396014 639390 396304 639406
rect 397670 639402 397960 639418
rect 397670 639396 397972 639402
rect 397670 639390 397920 639396
rect 386144 639338 386196 639344
rect 397920 639338 397972 639344
rect 398840 639396 398892 639402
rect 398840 639338 398892 639344
rect 370596 639328 370648 639334
rect 370596 639270 370648 639276
rect 370608 639268 370636 639270
rect 361488 639056 361540 639062
rect 361488 638998 361540 639004
rect 361212 598868 361264 598874
rect 361212 598810 361264 598816
rect 361120 598732 361172 598738
rect 361120 598674 361172 598680
rect 361028 598664 361080 598670
rect 361028 598606 361080 598612
rect 361040 553450 361068 598606
rect 361120 589960 361172 589966
rect 361120 589902 361172 589908
rect 361028 553444 361080 553450
rect 361028 553386 361080 553392
rect 360934 551984 360990 551993
rect 360934 551919 360990 551928
rect 361132 550662 361160 589902
rect 361500 552838 361528 638998
rect 398380 600296 398432 600302
rect 364550 600234 364840 600250
rect 398380 600238 398432 600244
rect 364550 600228 364852 600234
rect 364550 600222 364800 600228
rect 364800 600170 364852 600176
rect 365168 600228 365220 600234
rect 365168 600170 365220 600176
rect 361776 599078 361804 600100
rect 361868 600086 362342 600114
rect 361580 599072 361632 599078
rect 361580 599014 361632 599020
rect 361764 599072 361816 599078
rect 361764 599014 361816 599020
rect 361488 552832 361540 552838
rect 361488 552774 361540 552780
rect 361592 551857 361620 599014
rect 361868 586514 361896 600086
rect 362880 598176 362908 600100
rect 363248 600086 363446 600114
rect 362880 598148 363000 598176
rect 362972 595610 363000 598148
rect 362960 595604 363012 595610
rect 362960 595546 363012 595552
rect 361684 586486 361896 586514
rect 361684 560289 361712 586486
rect 363052 562420 363104 562426
rect 363052 562362 363104 562368
rect 361670 560280 361726 560289
rect 361670 560215 361726 560224
rect 362960 559700 363012 559706
rect 362960 559642 363012 559648
rect 361762 558920 361818 558929
rect 361762 558855 361818 558864
rect 361578 551848 361634 551857
rect 361578 551783 361634 551792
rect 361120 550656 361172 550662
rect 360842 550624 360898 550633
rect 361120 550598 361172 550604
rect 360842 550559 360898 550568
rect 361132 549930 361160 550598
rect 361776 549930 361804 558855
rect 362592 558272 362644 558278
rect 362592 558214 362644 558220
rect 362604 550118 362632 558214
rect 362972 550186 363000 559642
rect 363064 557534 363092 562362
rect 363064 557506 363184 557534
rect 362960 550180 363012 550186
rect 362960 550122 363012 550128
rect 362592 550112 362644 550118
rect 362592 550054 362644 550060
rect 361132 549902 361330 549930
rect 361776 549902 361974 549930
rect 362604 549916 362632 550054
rect 362972 549930 363000 550122
rect 363156 550066 363184 557506
rect 363248 551614 363276 600086
rect 363604 598596 363656 598602
rect 363604 598538 363656 598544
rect 363616 553489 363644 598538
rect 363984 596902 364012 600100
rect 364720 600086 365102 600114
rect 364432 598188 364484 598194
rect 364432 598130 364484 598136
rect 363972 596896 364024 596902
rect 363972 596838 364024 596844
rect 363602 553480 363658 553489
rect 363602 553415 363658 553424
rect 363236 551608 363288 551614
rect 363236 551550 363288 551556
rect 364444 550798 364472 598130
rect 364720 591394 364748 600086
rect 364708 591388 364760 591394
rect 364708 591330 364760 591336
rect 364524 552900 364576 552906
rect 364524 552842 364576 552848
rect 364432 550792 364484 550798
rect 364432 550734 364484 550740
rect 363156 550038 363552 550066
rect 363524 549930 363552 550038
rect 362972 549902 363262 549930
rect 363524 549902 363906 549930
rect 364536 549916 364564 552842
rect 365180 549930 365208 600170
rect 398392 600114 398420 600238
rect 365272 600086 365654 600114
rect 365272 598194 365300 600086
rect 365720 599616 365772 599622
rect 365720 599558 365772 599564
rect 365260 598188 365312 598194
rect 365260 598130 365312 598136
rect 364904 549916 365208 549930
rect 365732 549930 365760 599558
rect 366192 598534 366220 600100
rect 366284 600086 366758 600114
rect 366180 598528 366232 598534
rect 366180 598470 366232 598476
rect 366284 586514 366312 600086
rect 367296 598233 367324 600100
rect 367388 600086 367862 600114
rect 368032 600086 368414 600114
rect 368492 600086 368966 600114
rect 369044 600086 369518 600114
rect 369872 600086 370070 600114
rect 367282 598224 367338 598233
rect 367100 598188 367152 598194
rect 367282 598159 367338 598168
rect 367100 598130 367152 598136
rect 365824 586486 366312 586514
rect 365824 558890 365852 586486
rect 367112 567866 367140 598130
rect 367388 595542 367416 600086
rect 368032 598194 368060 600086
rect 368020 598188 368072 598194
rect 368020 598130 368072 598136
rect 367376 595536 367428 595542
rect 367376 595478 367428 595484
rect 367100 567860 367152 567866
rect 367100 567802 367152 567808
rect 365904 566500 365956 566506
rect 365904 566442 365956 566448
rect 365812 558884 365864 558890
rect 365812 558826 365864 558832
rect 365916 557534 365944 566442
rect 367376 565208 367428 565214
rect 367376 565150 367428 565156
rect 367192 563780 367244 563786
rect 367192 563722 367244 563728
rect 367204 557534 367232 563722
rect 367388 557534 367416 565150
rect 365916 557506 366128 557534
rect 367204 557506 367324 557534
rect 367388 557506 367968 557534
rect 366100 549930 366128 557506
rect 367100 552152 367152 552158
rect 367100 552094 367152 552100
rect 364904 549902 365194 549916
rect 365732 549902 365838 549930
rect 366100 549902 366482 549930
rect 367112 549916 367140 552094
rect 367296 549930 367324 557506
rect 367940 549930 367968 557506
rect 368492 554305 368520 600086
rect 369044 590034 369072 600086
rect 369032 590028 369084 590034
rect 369032 589970 369084 589976
rect 368572 584520 368624 584526
rect 368572 584462 368624 584468
rect 368584 557534 368612 584462
rect 368584 557506 369256 557534
rect 368478 554296 368534 554305
rect 368478 554231 368534 554240
rect 369030 552120 369086 552129
rect 369030 552055 369086 552064
rect 367296 549902 367770 549930
rect 367940 549902 368414 549930
rect 369044 549916 369072 552055
rect 369228 549930 369256 557506
rect 369872 554810 369900 600086
rect 370608 598369 370636 600100
rect 370594 598360 370650 598369
rect 370594 598295 370650 598304
rect 371160 598233 371188 600100
rect 371712 598602 371740 600100
rect 371804 600086 372278 600114
rect 372830 600086 372936 600114
rect 371700 598596 371752 598602
rect 371700 598538 371752 598544
rect 371146 598224 371202 598233
rect 371146 598159 371202 598168
rect 371804 588674 371832 600086
rect 372620 599684 372672 599690
rect 372620 599626 372672 599632
rect 371884 591388 371936 591394
rect 371884 591330 371936 591336
rect 371792 588668 371844 588674
rect 371792 588610 371844 588616
rect 369950 569256 370006 569265
rect 369950 569191 370006 569200
rect 369964 557534 369992 569191
rect 371608 558884 371660 558890
rect 371608 558826 371660 558832
rect 369964 557506 370544 557534
rect 369860 554804 369912 554810
rect 369860 554746 369912 554752
rect 369872 554130 369900 554746
rect 369860 554124 369912 554130
rect 369860 554066 369912 554072
rect 370516 549930 370544 557506
rect 371620 549930 371648 558826
rect 371896 552430 371924 591330
rect 371884 552424 371936 552430
rect 371884 552366 371936 552372
rect 369228 549902 369702 549930
rect 370516 549902 370990 549930
rect 371344 549916 371648 549930
rect 371896 549930 371924 552366
rect 372632 549930 372660 599626
rect 372804 598188 372856 598194
rect 372804 598130 372856 598136
rect 372712 598120 372764 598126
rect 372712 598062 372764 598068
rect 372724 557598 372752 598062
rect 372816 562426 372844 598130
rect 372908 587178 372936 600086
rect 373000 600086 373382 600114
rect 373552 600086 373934 600114
rect 374012 600086 374486 600114
rect 374564 600086 375038 600114
rect 375392 600086 375590 600114
rect 373000 598194 373028 600086
rect 372988 598188 373040 598194
rect 372988 598130 373040 598136
rect 373552 598126 373580 600086
rect 373540 598120 373592 598126
rect 373540 598062 373592 598068
rect 372896 587172 372948 587178
rect 372896 587114 372948 587120
rect 372804 562420 372856 562426
rect 372804 562362 372856 562368
rect 374012 558278 374040 600086
rect 374564 586514 374592 600086
rect 375392 594182 375420 600086
rect 376128 597689 376156 600100
rect 376680 598194 376708 600100
rect 377232 598602 377260 600100
rect 377324 600086 377798 600114
rect 378244 600086 378350 600114
rect 377220 598596 377272 598602
rect 377220 598538 377272 598544
rect 376668 598188 376720 598194
rect 376668 598130 376720 598136
rect 376114 597680 376170 597689
rect 376114 597615 376170 597624
rect 375380 594176 375432 594182
rect 375380 594118 375432 594124
rect 377324 586514 377352 600086
rect 377404 598188 377456 598194
rect 377404 598130 377456 598136
rect 374104 586486 374592 586514
rect 376772 586486 377352 586514
rect 374104 559706 374132 586486
rect 374276 580304 374328 580310
rect 374276 580246 374328 580252
rect 374092 559700 374144 559706
rect 374092 559642 374144 559648
rect 374000 558272 374052 558278
rect 374000 558214 374052 558220
rect 372712 557592 372764 557598
rect 372712 557534 372764 557540
rect 374288 557534 374316 580246
rect 376772 576881 376800 586486
rect 376758 576872 376814 576881
rect 376758 576807 376814 576816
rect 376944 573436 376996 573442
rect 376944 573378 376996 573384
rect 375380 562352 375432 562358
rect 375380 562294 375432 562300
rect 372724 557054 372752 557534
rect 374288 557506 374408 557534
rect 372712 557048 372764 557054
rect 372712 556990 372764 556996
rect 374184 552832 374236 552838
rect 374184 552774 374236 552780
rect 373540 552084 373592 552090
rect 373540 552026 373592 552032
rect 371344 549902 371634 549916
rect 371896 549902 372278 549930
rect 372632 549902 372922 549930
rect 373552 549916 373580 552026
rect 374196 549916 374224 552774
rect 374380 549930 374408 557506
rect 375392 549930 375420 562294
rect 376852 558272 376904 558278
rect 376852 558214 376904 558220
rect 376864 553382 376892 558214
rect 376852 553376 376904 553382
rect 376852 553318 376904 553324
rect 376760 553036 376812 553042
rect 376760 552978 376812 552984
rect 376116 552832 376168 552838
rect 376116 552774 376168 552780
rect 374380 549902 374854 549930
rect 375392 549902 375498 549930
rect 376128 549916 376156 552774
rect 376772 549916 376800 552978
rect 376956 549930 376984 573378
rect 377416 551070 377444 598130
rect 378244 563961 378272 600086
rect 378416 599752 378468 599758
rect 378416 599694 378468 599700
rect 378324 598188 378376 598194
rect 378324 598130 378376 598136
rect 378336 583137 378364 598130
rect 378322 583128 378378 583137
rect 378322 583063 378378 583072
rect 378230 563952 378286 563961
rect 378230 563887 378286 563896
rect 378428 557534 378456 599694
rect 378888 598233 378916 600100
rect 379072 600086 379454 600114
rect 379716 600086 380006 600114
rect 380176 600086 380558 600114
rect 378874 598224 378930 598233
rect 379072 598194 379100 600086
rect 378874 598159 378930 598168
rect 379060 598188 379112 598194
rect 379060 598130 379112 598136
rect 379612 598188 379664 598194
rect 379612 598130 379664 598136
rect 378428 557506 379008 557534
rect 377772 553376 377824 553382
rect 377772 553318 377824 553324
rect 377404 551064 377456 551070
rect 377404 551006 377456 551012
rect 377784 549930 377812 553318
rect 378692 553104 378744 553110
rect 378692 553046 378744 553052
rect 377956 551064 378008 551070
rect 377956 551006 378008 551012
rect 377968 550050 377996 551006
rect 377956 550044 378008 550050
rect 377956 549986 378008 549992
rect 376956 549902 377430 549930
rect 377784 549902 378074 549930
rect 378704 549916 378732 553046
rect 378980 549930 379008 557506
rect 379624 556918 379652 598130
rect 379716 581913 379744 600086
rect 379796 599820 379848 599826
rect 379796 599762 379848 599768
rect 379702 581904 379758 581913
rect 379702 581839 379758 581848
rect 379612 556912 379664 556918
rect 379612 556854 379664 556860
rect 379808 549930 379836 599762
rect 380176 598194 380204 600086
rect 381096 598670 381124 600100
rect 381188 600086 381662 600114
rect 381832 600086 382214 600114
rect 382476 600086 382766 600114
rect 382936 600086 383318 600114
rect 383672 600086 383870 600114
rect 381084 598664 381136 598670
rect 381084 598606 381136 598612
rect 380164 598188 380216 598194
rect 380164 598130 380216 598136
rect 380992 598188 381044 598194
rect 380992 598130 381044 598136
rect 381004 563718 381032 598130
rect 381084 565140 381136 565146
rect 381084 565082 381136 565088
rect 380992 563712 381044 563718
rect 380992 563654 381044 563660
rect 380624 552764 380676 552770
rect 380624 552706 380676 552712
rect 378980 549902 379362 549930
rect 379808 549902 380006 549930
rect 380636 549916 380664 552706
rect 381096 549930 381124 565082
rect 381188 558346 381216 600086
rect 381832 598194 381860 600086
rect 382280 599888 382332 599894
rect 382280 599830 382332 599836
rect 381820 598188 381872 598194
rect 381820 598130 381872 598136
rect 381544 594176 381596 594182
rect 381544 594118 381596 594124
rect 381176 558340 381228 558346
rect 381176 558282 381228 558288
rect 381556 552362 381584 594118
rect 381544 552356 381596 552362
rect 381544 552298 381596 552304
rect 381556 549930 381584 552298
rect 382292 551274 382320 599830
rect 382372 598188 382424 598194
rect 382372 598130 382424 598136
rect 382384 565185 382412 598130
rect 382476 581777 382504 600086
rect 382936 598194 382964 600086
rect 382924 598188 382976 598194
rect 382924 598130 382976 598136
rect 382462 581768 382518 581777
rect 382462 581703 382518 581712
rect 382464 574796 382516 574802
rect 382464 574738 382516 574744
rect 382370 565176 382426 565185
rect 382370 565111 382426 565120
rect 382280 551268 382332 551274
rect 382280 551210 382332 551216
rect 382476 549930 382504 574738
rect 383672 551682 383700 600086
rect 384408 596630 384436 600100
rect 384500 600086 384974 600114
rect 385144 600086 385526 600114
rect 385696 600086 386078 600114
rect 386524 600086 386630 600114
rect 384396 596624 384448 596630
rect 384396 596566 384448 596572
rect 384500 586514 384528 600086
rect 385040 598188 385092 598194
rect 385040 598130 385092 598136
rect 383764 586486 384528 586514
rect 383764 552770 383792 586486
rect 383844 562420 383896 562426
rect 383844 562362 383896 562368
rect 383752 552764 383804 552770
rect 383752 552706 383804 552712
rect 383660 551676 383712 551682
rect 383660 551618 383712 551624
rect 382924 551268 382976 551274
rect 382924 551210 382976 551216
rect 382936 549930 382964 551210
rect 383856 549930 383884 562362
rect 385052 555558 385080 598130
rect 385144 565554 385172 600086
rect 385696 598194 385724 600086
rect 386420 598868 386472 598874
rect 386420 598810 386472 598816
rect 385684 598188 385736 598194
rect 385684 598130 385736 598136
rect 386432 594182 386460 598810
rect 386420 594176 386472 594182
rect 386420 594118 386472 594124
rect 385684 589280 385736 589286
rect 385684 589222 385736 589228
rect 385132 565548 385184 565554
rect 385132 565490 385184 565496
rect 385040 555552 385092 555558
rect 385040 555494 385092 555500
rect 385696 552226 385724 589222
rect 385776 582412 385828 582418
rect 385776 582354 385828 582360
rect 385788 552430 385816 582354
rect 386524 559638 386552 600086
rect 386604 599004 386656 599010
rect 386604 598946 386656 598952
rect 386616 580417 386644 598946
rect 387168 598874 387196 600100
rect 387720 599146 387748 600100
rect 387708 599140 387760 599146
rect 387708 599082 387760 599088
rect 387720 599010 387748 599082
rect 387708 599004 387760 599010
rect 387708 598946 387760 598952
rect 388272 598942 388300 600100
rect 388456 600086 388838 600114
rect 389192 600086 389390 600114
rect 389560 600086 389942 600114
rect 390112 600086 390494 600114
rect 390664 600086 391046 600114
rect 391216 600086 391598 600114
rect 391952 600086 392150 600114
rect 392228 600086 392702 600114
rect 392780 600086 393254 600114
rect 393424 600086 393806 600114
rect 393976 600086 394358 600114
rect 394804 600086 394910 600114
rect 395080 600086 395462 600114
rect 395540 600086 396014 600114
rect 396184 600086 396566 600114
rect 396736 600086 397118 600114
rect 397564 600086 397670 600114
rect 398222 600100 398420 600114
rect 398208 600086 398420 600100
rect 388260 598936 388312 598942
rect 388260 598878 388312 598884
rect 387156 598868 387208 598874
rect 387156 598810 387208 598816
rect 388272 598194 388300 598878
rect 388456 598806 388484 600086
rect 388444 598800 388496 598806
rect 388444 598742 388496 598748
rect 388260 598188 388312 598194
rect 388260 598130 388312 598136
rect 387800 595604 387852 595610
rect 387800 595546 387852 595552
rect 386788 591320 386840 591326
rect 386788 591262 386840 591268
rect 386602 580408 386658 580417
rect 386602 580343 386658 580352
rect 386604 576156 386656 576162
rect 386604 576098 386656 576104
rect 386512 559632 386564 559638
rect 386512 559574 386564 559580
rect 385776 552424 385828 552430
rect 385776 552366 385828 552372
rect 384488 552220 384540 552226
rect 384488 552162 384540 552168
rect 385684 552220 385736 552226
rect 385684 552162 385736 552168
rect 384500 551002 384528 552162
rect 384488 550996 384540 551002
rect 384488 550938 384540 550944
rect 381096 549902 381294 549930
rect 381556 549902 381938 549930
rect 382476 549902 382582 549930
rect 382936 549902 383226 549930
rect 383672 549916 383884 549930
rect 384500 549916 384528 550938
rect 385788 549916 385816 552366
rect 386616 550322 386644 576098
rect 386696 560992 386748 560998
rect 386696 560934 386748 560940
rect 386708 550634 386736 560934
rect 386800 557534 386828 591262
rect 387812 576854 387840 595546
rect 387812 576826 387932 576854
rect 387904 557534 387932 576826
rect 388456 560289 388484 598742
rect 388536 598188 388588 598194
rect 388536 598130 388588 598136
rect 388548 568041 388576 598130
rect 388628 568608 388680 568614
rect 388628 568550 388680 568556
rect 388534 568032 388590 568041
rect 388534 567967 388590 567976
rect 388442 560280 388498 560289
rect 388442 560215 388498 560224
rect 386800 557506 387288 557534
rect 387904 557506 388024 557534
rect 386708 550606 386828 550634
rect 386604 550316 386656 550322
rect 386604 550258 386656 550264
rect 386800 549930 386828 550606
rect 387064 550316 387116 550322
rect 387064 550258 387116 550264
rect 383672 549902 383870 549916
rect 386446 549902 386828 549930
rect 387076 549916 387104 550258
rect 387260 549930 387288 557506
rect 387996 552362 388024 557506
rect 387984 552356 388036 552362
rect 387984 552298 388036 552304
rect 387996 549930 388024 552298
rect 388640 551138 388668 568550
rect 389192 551750 389220 600086
rect 389272 598188 389324 598194
rect 389272 598130 389324 598136
rect 389284 582418 389312 598130
rect 389560 586514 389588 600086
rect 390112 598194 390140 600086
rect 390100 598188 390152 598194
rect 390100 598130 390152 598136
rect 390560 597644 390612 597650
rect 390560 597586 390612 597592
rect 389376 586486 389588 586514
rect 389376 583817 389404 586486
rect 389362 583808 389418 583817
rect 389362 583743 389418 583752
rect 389272 582412 389324 582418
rect 389272 582354 389324 582360
rect 389272 572008 389324 572014
rect 389272 571950 389324 571956
rect 389284 557534 389312 571950
rect 390572 562494 390600 597586
rect 390664 589286 390692 600086
rect 391216 597650 391244 600086
rect 391204 597644 391256 597650
rect 391204 597586 391256 597592
rect 391202 596864 391258 596873
rect 391202 596799 391258 596808
rect 390652 589280 390704 589286
rect 390652 589222 390704 589228
rect 390652 576224 390704 576230
rect 390652 576166 390704 576172
rect 390560 562488 390612 562494
rect 390560 562430 390612 562436
rect 389284 557506 389864 557534
rect 389640 552900 389692 552906
rect 389640 552842 389692 552848
rect 389180 551744 389232 551750
rect 389180 551686 389232 551692
rect 388628 551132 388680 551138
rect 388628 551074 388680 551080
rect 388996 551132 389048 551138
rect 388996 551074 389048 551080
rect 387260 549902 387734 549930
rect 387996 549902 388378 549930
rect 389008 549916 389036 551074
rect 389652 549916 389680 552842
rect 389836 549930 389864 557506
rect 390664 549930 390692 576166
rect 391216 550662 391244 596799
rect 391952 589966 391980 600086
rect 392228 598210 392256 600086
rect 392044 598182 392256 598210
rect 392044 591394 392072 598182
rect 392780 596714 392808 600086
rect 393320 598188 393372 598194
rect 393320 598130 393372 598136
rect 392136 596686 392808 596714
rect 392136 595513 392164 596686
rect 392584 596624 392636 596630
rect 392584 596566 392636 596572
rect 392122 595504 392178 595513
rect 392122 595439 392178 595448
rect 392032 591388 392084 591394
rect 392032 591330 392084 591336
rect 391940 589960 391992 589966
rect 391940 589902 391992 589908
rect 391940 565548 391992 565554
rect 391940 565490 391992 565496
rect 391204 550656 391256 550662
rect 391204 550598 391256 550604
rect 391216 549930 391244 550598
rect 391952 549930 391980 565490
rect 392596 553382 392624 596566
rect 392584 553376 392636 553382
rect 392584 553318 392636 553324
rect 392860 553036 392912 553042
rect 392860 552978 392912 552984
rect 389836 549902 390310 549930
rect 390664 549902 390954 549930
rect 391216 549902 391598 549930
rect 391952 549902 392242 549930
rect 392872 549916 392900 552978
rect 393332 552022 393360 598130
rect 393424 568614 393452 600086
rect 393976 598194 394004 600086
rect 393964 598188 394016 598194
rect 393964 598130 394016 598136
rect 394700 598188 394752 598194
rect 394700 598130 394752 598136
rect 393412 568608 393464 568614
rect 393412 568550 393464 568556
rect 394148 553376 394200 553382
rect 394148 553318 394200 553324
rect 393504 552492 393556 552498
rect 393504 552434 393556 552440
rect 393320 552016 393372 552022
rect 393320 551958 393372 551964
rect 393516 549916 393544 552434
rect 394160 549916 394188 553318
rect 394712 550050 394740 598130
rect 394804 566574 394832 600086
rect 395080 598194 395108 600086
rect 395068 598188 395120 598194
rect 395068 598130 395120 598136
rect 395540 586673 395568 600086
rect 396080 598188 396132 598194
rect 396080 598130 396132 598136
rect 395526 586664 395582 586673
rect 395526 586599 395582 586608
rect 394884 570648 394936 570654
rect 394884 570590 394936 570596
rect 394792 566568 394844 566574
rect 394792 566510 394844 566516
rect 394896 557534 394924 570590
rect 394896 557506 395016 557534
rect 394792 552220 394844 552226
rect 394792 552162 394844 552168
rect 394700 550044 394752 550050
rect 394700 549986 394752 549992
rect 394804 549916 394832 552162
rect 394988 549930 395016 557506
rect 396092 556850 396120 598130
rect 396184 584594 396212 600086
rect 396736 598194 396764 600086
rect 396724 598188 396776 598194
rect 396724 598130 396776 598136
rect 396722 585712 396778 585721
rect 396722 585647 396778 585656
rect 396172 584588 396224 584594
rect 396172 584530 396224 584536
rect 396080 556844 396132 556850
rect 396080 556786 396132 556792
rect 396356 552968 396408 552974
rect 396356 552910 396408 552916
rect 396080 550792 396132 550798
rect 396080 550734 396132 550740
rect 394988 549902 395462 549930
rect 396092 549916 396120 550734
rect 396368 549930 396396 552910
rect 396736 552294 396764 585647
rect 397368 552696 397420 552702
rect 397368 552638 397420 552644
rect 396724 552288 396776 552294
rect 396724 552230 396776 552236
rect 396368 549902 396750 549930
rect 397380 549916 397408 552638
rect 397460 550928 397512 550934
rect 397460 550870 397512 550876
rect 397472 550633 397500 550870
rect 397458 550624 397514 550633
rect 397458 550559 397514 550568
rect 397564 550526 397592 600086
rect 397644 598596 397696 598602
rect 397644 598538 397696 598544
rect 397552 550520 397604 550526
rect 397552 550462 397604 550468
rect 397656 549914 397684 598538
rect 397736 598528 397788 598534
rect 397736 598470 397788 598476
rect 397748 576854 397776 598470
rect 398208 596834 398236 600086
rect 398196 596828 398248 596834
rect 398196 596770 398248 596776
rect 397748 576826 398144 576854
rect 398012 552288 398064 552294
rect 398012 552230 398064 552236
rect 398024 549916 398052 552230
rect 398116 550633 398144 576826
rect 398656 552288 398708 552294
rect 398656 552230 398708 552236
rect 398102 550624 398158 550633
rect 398102 550559 398158 550568
rect 398668 549916 398696 552230
rect 398852 549930 398880 639338
rect 398944 553042 398972 639934
rect 399024 639464 399076 639470
rect 399024 639406 399076 639412
rect 398932 553036 398984 553042
rect 398932 552978 398984 552984
rect 399036 552838 399064 639406
rect 399024 552832 399076 552838
rect 399024 552774 399076 552780
rect 399128 552498 399156 642398
rect 399208 642388 399260 642394
rect 399208 642330 399260 642336
rect 399220 599826 399248 642330
rect 399208 599820 399260 599826
rect 399208 599762 399260 599768
rect 399312 599758 399340 642602
rect 400312 642592 400364 642598
rect 400312 642534 400364 642540
rect 399668 642116 399720 642122
rect 399668 642058 399720 642064
rect 399392 641844 399444 641850
rect 399392 641786 399444 641792
rect 399300 599752 399352 599758
rect 399300 599694 399352 599700
rect 399404 599690 399432 641786
rect 399392 599684 399444 599690
rect 399392 599626 399444 599632
rect 399574 559600 399630 559609
rect 399574 559535 399630 559544
rect 399484 552764 399536 552770
rect 399484 552706 399536 552712
rect 399116 552492 399168 552498
rect 399116 552434 399168 552440
rect 397644 549908 397696 549914
rect 364904 549846 364932 549902
rect 371344 549846 371372 549902
rect 383672 549846 383700 549902
rect 398852 549902 399326 549930
rect 397644 549850 397696 549856
rect 364892 549840 364944 549846
rect 364892 549782 364944 549788
rect 371332 549840 371384 549846
rect 371332 549782 371384 549788
rect 383660 549840 383712 549846
rect 383660 549782 383712 549788
rect 359568 538186 359780 538214
rect 359464 530324 359516 530330
rect 359464 530266 359516 530272
rect 359568 529666 359596 538186
rect 359740 534132 359792 534138
rect 359740 534074 359792 534080
rect 359752 529904 359780 534074
rect 359832 530052 359884 530058
rect 359884 530000 359964 530006
rect 359832 529994 359964 530000
rect 359844 529978 359964 529994
rect 359752 529876 359872 529904
rect 359568 529638 359780 529666
rect 359370 528320 359426 528329
rect 359370 528255 359426 528264
rect 359648 522980 359700 522986
rect 359648 522922 359700 522928
rect 359278 520976 359334 520985
rect 359278 520911 359334 520920
rect 359556 514888 359608 514894
rect 359556 514830 359608 514836
rect 359002 513360 359058 513369
rect 359002 513295 359058 513304
rect 359464 513324 359516 513330
rect 359464 513266 359516 513272
rect 359372 500812 359424 500818
rect 359372 500754 359424 500760
rect 359384 497418 359412 500754
rect 359372 497412 359424 497418
rect 359372 497354 359424 497360
rect 358912 489184 358964 489190
rect 358912 489126 358964 489132
rect 358820 86964 358872 86970
rect 358820 86906 358872 86912
rect 359476 6866 359504 513266
rect 359568 46918 359596 514830
rect 359660 245614 359688 522922
rect 359752 507890 359780 529638
rect 359740 507884 359792 507890
rect 359740 507826 359792 507832
rect 359740 505164 359792 505170
rect 359740 505106 359792 505112
rect 359752 499186 359780 505106
rect 359844 499254 359872 529876
rect 359832 499248 359884 499254
rect 359832 499190 359884 499196
rect 359740 499180 359792 499186
rect 359740 499122 359792 499128
rect 359936 499118 359964 529978
rect 399496 507385 399524 552706
rect 399588 523705 399616 559535
rect 399680 525774 399708 642058
rect 399760 641776 399812 641782
rect 399760 641718 399812 641724
rect 399772 550594 399800 641718
rect 400220 639328 400272 639334
rect 400220 639270 400272 639276
rect 399944 561060 399996 561066
rect 399944 561002 399996 561008
rect 399852 551744 399904 551750
rect 399852 551686 399904 551692
rect 399760 550588 399812 550594
rect 399760 550530 399812 550536
rect 399864 536625 399892 551686
rect 399956 546145 399984 561002
rect 400036 551676 400088 551682
rect 400036 551618 400088 551624
rect 399942 546136 399998 546145
rect 399942 546071 399998 546080
rect 400048 541566 400076 551618
rect 400126 541580 400182 541589
rect 400048 541538 400126 541566
rect 400126 541515 400182 541524
rect 399850 536616 399906 536625
rect 399850 536551 399906 536560
rect 399758 535664 399814 535673
rect 399758 535599 399814 535608
rect 399772 533225 399800 535599
rect 399758 533216 399814 533225
rect 399758 533151 399814 533160
rect 399668 525768 399720 525774
rect 399668 525710 399720 525716
rect 399574 523696 399630 523705
rect 399574 523631 399630 523640
rect 399482 507376 399538 507385
rect 399482 507311 399538 507320
rect 400232 504189 400260 639270
rect 400324 525269 400352 642534
rect 403164 642524 403216 642530
rect 403164 642466 403216 642472
rect 400496 642320 400548 642326
rect 400496 642262 400548 642268
rect 400862 642288 400918 642297
rect 400404 639124 400456 639130
rect 400404 639066 400456 639072
rect 400416 552906 400444 639066
rect 400508 599622 400536 642262
rect 400862 642223 400918 642232
rect 400956 642252 401008 642258
rect 400588 641912 400640 641918
rect 400588 641854 400640 641860
rect 400600 599894 400628 641854
rect 400588 599888 400640 599894
rect 400588 599830 400640 599836
rect 400496 599616 400548 599622
rect 400496 599558 400548 599564
rect 400494 561096 400550 561105
rect 400494 561031 400550 561040
rect 400404 552900 400456 552906
rect 400404 552842 400456 552848
rect 400404 551608 400456 551614
rect 400404 551550 400456 551556
rect 400416 535469 400444 551550
rect 400402 535460 400458 535469
rect 400402 535395 400458 535404
rect 400310 525260 400366 525269
rect 400310 525195 400366 525204
rect 400508 523025 400536 561031
rect 400588 552016 400640 552022
rect 400588 551958 400640 551964
rect 400494 523016 400550 523025
rect 400494 522951 400550 522960
rect 400600 515545 400628 551958
rect 400680 550520 400732 550526
rect 400680 550462 400732 550468
rect 400692 527105 400720 550462
rect 400772 550044 400824 550050
rect 400772 549986 400824 549992
rect 400784 538121 400812 549986
rect 400770 538112 400826 538121
rect 400770 538047 400826 538056
rect 400770 536344 400826 536353
rect 400770 536279 400826 536288
rect 400678 527096 400734 527105
rect 400678 527031 400734 527040
rect 400586 515536 400642 515545
rect 400586 515471 400642 515480
rect 400218 504180 400274 504189
rect 400218 504115 400274 504124
rect 399482 501664 399538 501673
rect 399482 501599 399538 501608
rect 399496 500954 399524 501599
rect 399484 500948 399536 500954
rect 399484 500890 399536 500896
rect 359924 499112 359976 499118
rect 359924 499054 359976 499060
rect 360028 498137 360056 500140
rect 360672 499905 360700 500140
rect 360844 499996 360896 500002
rect 360844 499938 360896 499944
rect 360658 499896 360714 499905
rect 360658 499831 360714 499840
rect 360014 498128 360070 498137
rect 360014 498063 360070 498072
rect 360856 497185 360884 499938
rect 361316 498166 361344 500140
rect 361960 499225 361988 500140
rect 362604 499905 362632 500140
rect 362590 499896 362646 499905
rect 362590 499831 362646 499840
rect 361946 499216 362002 499225
rect 361946 499151 362002 499160
rect 362960 498840 363012 498846
rect 362960 498782 363012 498788
rect 361304 498160 361356 498166
rect 361304 498102 361356 498108
rect 362972 497729 363000 498782
rect 363248 497758 363276 500140
rect 363892 497865 363920 500140
rect 364536 499526 364564 500140
rect 365180 499905 365208 500140
rect 365166 499896 365222 499905
rect 365166 499831 365222 499840
rect 364524 499520 364576 499526
rect 365824 499497 365852 500140
rect 364524 499462 364576 499468
rect 365810 499488 365866 499497
rect 365810 499423 365866 499432
rect 363878 497856 363934 497865
rect 363878 497791 363934 497800
rect 364062 497856 364118 497865
rect 366468 497826 366496 500140
rect 367112 498030 367140 500140
rect 367756 499497 367784 500140
rect 368400 499905 368428 500140
rect 368386 499896 368442 499905
rect 368386 499831 368442 499840
rect 367742 499488 367798 499497
rect 367742 499423 367798 499432
rect 367756 498914 367784 499423
rect 367744 498908 367796 498914
rect 367744 498850 367796 498856
rect 367100 498024 367152 498030
rect 369044 498001 369072 500140
rect 369688 499905 369716 500140
rect 370332 499905 370360 500140
rect 369674 499896 369730 499905
rect 369674 499831 369730 499840
rect 370318 499896 370374 499905
rect 370318 499831 370374 499840
rect 370976 498098 371004 500140
rect 371620 498953 371648 500140
rect 371606 498944 371662 498953
rect 371606 498879 371662 498888
rect 370964 498092 371016 498098
rect 370964 498034 371016 498040
rect 367100 497966 367152 497972
rect 369030 497992 369086 498001
rect 369030 497927 369086 497936
rect 364062 497791 364118 497800
rect 366456 497820 366508 497826
rect 363236 497752 363288 497758
rect 362958 497720 363014 497729
rect 363236 497694 363288 497700
rect 362958 497655 363014 497664
rect 364076 497457 364104 497791
rect 366456 497762 366508 497768
rect 372264 497622 372292 500140
rect 372252 497616 372304 497622
rect 372252 497558 372304 497564
rect 364062 497448 364118 497457
rect 364062 497383 364118 497392
rect 360842 497176 360898 497185
rect 360842 497111 360898 497120
rect 366364 496800 366416 496806
rect 366364 496742 366416 496748
rect 362224 494012 362276 494018
rect 362224 493954 362276 493960
rect 362236 353258 362264 493954
rect 364340 482316 364392 482322
rect 364340 482258 364392 482264
rect 362224 353252 362276 353258
rect 362224 353194 362276 353200
rect 359648 245608 359700 245614
rect 359648 245550 359700 245556
rect 359556 46912 359608 46918
rect 359556 46854 359608 46860
rect 360200 18760 360252 18766
rect 360200 18702 360252 18708
rect 360212 16574 360240 18702
rect 364352 16574 364380 482258
rect 366376 405686 366404 496742
rect 367100 496120 367152 496126
rect 367100 496062 367152 496068
rect 366364 405680 366416 405686
rect 366364 405622 366416 405628
rect 367112 16574 367140 496062
rect 369124 494760 369176 494766
rect 369124 494702 369176 494708
rect 369136 59362 369164 494702
rect 372908 126954 372936 500140
rect 373552 499458 373580 500140
rect 374840 499905 374868 500140
rect 374826 499896 374882 499905
rect 374826 499831 374882 499840
rect 373540 499452 373592 499458
rect 373540 499394 373592 499400
rect 375484 498710 375512 500140
rect 376128 499905 376156 500140
rect 376772 499905 376800 500140
rect 376114 499896 376170 499905
rect 376114 499831 376170 499840
rect 376758 499896 376814 499905
rect 376758 499831 376814 499840
rect 375472 498704 375524 498710
rect 375472 498646 375524 498652
rect 376128 497457 376156 499831
rect 377416 499497 377444 500140
rect 377402 499488 377458 499497
rect 377402 499423 377458 499432
rect 378060 498642 378088 500140
rect 378048 498636 378100 498642
rect 378048 498578 378100 498584
rect 376114 497448 376170 497457
rect 376114 497383 376170 497392
rect 374000 479528 374052 479534
rect 374000 479470 374052 479476
rect 372896 126948 372948 126954
rect 372896 126890 372948 126896
rect 369124 59356 369176 59362
rect 369124 59298 369176 59304
rect 371240 22772 371292 22778
rect 371240 22714 371292 22720
rect 360212 16546 361160 16574
rect 364352 16546 364656 16574
rect 367112 16546 367784 16574
rect 359464 6860 359516 6866
rect 359464 6802 359516 6808
rect 357624 5024 357676 5030
rect 357624 4966 357676 4972
rect 361132 480 361160 16546
rect 364628 480 364656 16546
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 22714
rect 374012 3058 374040 479470
rect 378140 31068 378192 31074
rect 378140 31010 378192 31016
rect 378152 16574 378180 31010
rect 378152 16546 378456 16574
rect 374000 3052 374052 3058
rect 374000 2994 374052 3000
rect 375288 3052 375340 3058
rect 375288 2994 375340 3000
rect 375300 480 375328 2994
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378704 11762 378732 500140
rect 379348 497962 379376 500140
rect 379336 497956 379388 497962
rect 379336 497898 379388 497904
rect 379992 497894 380020 500140
rect 380636 499905 380664 500140
rect 381280 499905 381308 500140
rect 380622 499896 380678 499905
rect 380622 499831 380678 499840
rect 381266 499896 381322 499905
rect 381266 499831 381322 499840
rect 381924 498982 381952 500140
rect 382568 499905 382596 500140
rect 382554 499896 382610 499905
rect 382554 499831 382610 499840
rect 381912 498976 381964 498982
rect 381912 498918 381964 498924
rect 379980 497888 380032 497894
rect 379980 497830 380032 497836
rect 382568 497593 382596 499831
rect 382554 497584 382610 497593
rect 382554 497519 382610 497528
rect 381544 496868 381596 496874
rect 381544 496810 381596 496816
rect 381556 225826 381584 496810
rect 382280 480956 382332 480962
rect 382280 480898 382332 480904
rect 381544 225820 381596 225826
rect 381544 225762 381596 225768
rect 382292 16574 382320 480898
rect 383212 299470 383240 500140
rect 383856 497350 383884 500140
rect 383844 497344 383896 497350
rect 383844 497286 383896 497292
rect 384500 496874 384528 500140
rect 385144 499905 385172 500140
rect 385130 499896 385186 499905
rect 385130 499831 385186 499840
rect 385144 497865 385172 499831
rect 385130 497856 385186 497865
rect 385130 497791 385186 497800
rect 385788 497729 385816 500140
rect 385774 497720 385830 497729
rect 385774 497655 385830 497664
rect 386432 497321 386460 500140
rect 387076 498137 387104 500140
rect 387062 498128 387118 498137
rect 387062 498063 387118 498072
rect 387720 498001 387748 500140
rect 388364 498030 388392 500140
rect 389652 498778 389680 500140
rect 390296 499905 390324 500140
rect 390282 499896 390338 499905
rect 390282 499831 390338 499840
rect 389640 498772 389692 498778
rect 389640 498714 389692 498720
rect 388352 498024 388404 498030
rect 387706 497992 387762 498001
rect 388352 497966 388404 497972
rect 387706 497927 387762 497936
rect 386418 497312 386474 497321
rect 386418 497247 386474 497256
rect 384488 496868 384540 496874
rect 384488 496810 384540 496816
rect 389180 493332 389232 493338
rect 389180 493274 389232 493280
rect 385040 478168 385092 478174
rect 385040 478110 385092 478116
rect 383200 299464 383252 299470
rect 383200 299406 383252 299412
rect 385052 16574 385080 478110
rect 389192 16574 389220 493274
rect 382292 16546 382412 16574
rect 385052 16546 386000 16574
rect 389192 16546 389496 16574
rect 378692 11756 378744 11762
rect 378692 11698 378744 11704
rect 382384 480 382412 16546
rect 385972 480 386000 16546
rect 389468 480 389496 16546
rect 390940 15978 390968 500140
rect 391584 499769 391612 500140
rect 391570 499760 391626 499769
rect 391570 499695 391626 499704
rect 391584 497185 391612 499695
rect 391570 497176 391626 497185
rect 391570 497111 391626 497120
rect 392228 491978 392256 500140
rect 392872 499905 392900 500140
rect 392858 499896 392914 499905
rect 392858 499831 392914 499840
rect 393516 499633 393544 500140
rect 393502 499624 393558 499633
rect 393502 499559 393558 499568
rect 394160 499526 394188 500140
rect 394148 499520 394200 499526
rect 394148 499462 394200 499468
rect 394804 497690 394832 500140
rect 395448 498137 395476 500140
rect 395434 498128 395490 498137
rect 395434 498063 395490 498072
rect 394792 497684 394844 497690
rect 394792 497626 394844 497632
rect 392216 491972 392268 491978
rect 392216 491914 392268 491920
rect 391940 476808 391992 476814
rect 391940 476750 391992 476756
rect 391952 16574 391980 476750
rect 391952 16546 392624 16574
rect 390928 15972 390980 15978
rect 390928 15914 390980 15920
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 396092 8294 396120 500140
rect 396736 498098 396764 500140
rect 397380 499050 397408 500140
rect 398024 499322 398052 500140
rect 398668 499905 398696 500140
rect 398654 499896 398710 499905
rect 398654 499831 398710 499840
rect 398012 499316 398064 499322
rect 398012 499258 398064 499264
rect 397368 499044 397420 499050
rect 397368 498986 397420 498992
rect 399312 498166 399340 500140
rect 400784 499390 400812 536279
rect 400876 529990 400904 642223
rect 400956 642194 401008 642200
rect 400968 540705 400996 642194
rect 401876 640688 401928 640694
rect 401876 640630 401928 640636
rect 401600 640620 401652 640626
rect 401600 640562 401652 640568
rect 401048 598460 401100 598466
rect 401048 598402 401100 598408
rect 400954 540696 401010 540705
rect 400954 540631 401010 540640
rect 401060 539345 401088 598402
rect 401612 547505 401640 640562
rect 401784 639600 401836 639606
rect 401784 639542 401836 639548
rect 401690 551576 401746 551585
rect 401690 551511 401746 551520
rect 401598 547496 401654 547505
rect 401598 547431 401654 547440
rect 401704 544785 401732 551511
rect 401690 544776 401746 544785
rect 401690 544711 401746 544720
rect 401600 543448 401652 543454
rect 401600 543390 401652 543396
rect 401612 543153 401640 543390
rect 401598 543144 401654 543153
rect 401598 543079 401654 543088
rect 401598 541784 401654 541793
rect 401598 541719 401654 541728
rect 401612 541006 401640 541719
rect 401600 541000 401652 541006
rect 401600 540942 401652 540948
rect 401046 539336 401102 539345
rect 401046 539271 401102 539280
rect 401600 536240 401652 536246
rect 401598 536208 401600 536217
rect 401652 536208 401654 536217
rect 401598 536143 401654 536152
rect 401796 533225 401824 639542
rect 401888 534721 401916 640630
rect 402336 639260 402388 639266
rect 402336 639202 402388 639208
rect 401968 639192 402020 639198
rect 401968 639134 402020 639140
rect 401980 540977 402008 639134
rect 402152 561128 402204 561134
rect 402152 561070 402204 561076
rect 402060 550588 402112 550594
rect 402060 550530 402112 550536
rect 401966 540968 402022 540977
rect 401966 540903 402022 540912
rect 401874 534712 401930 534721
rect 401874 534647 401930 534656
rect 401876 533792 401928 533798
rect 401874 533760 401876 533769
rect 401928 533760 401930 533769
rect 401874 533695 401930 533704
rect 401782 533216 401838 533225
rect 401782 533151 401838 533160
rect 401968 531956 402020 531962
rect 401968 531898 402020 531904
rect 401980 531865 402008 531898
rect 401966 531856 402022 531865
rect 401966 531791 402022 531800
rect 401968 531276 402020 531282
rect 401968 531218 402020 531224
rect 401980 530233 402008 531218
rect 401966 530224 402022 530233
rect 401966 530159 402022 530168
rect 400864 529984 400916 529990
rect 400864 529926 400916 529932
rect 401876 529984 401928 529990
rect 401876 529926 401928 529932
rect 401782 527096 401838 527105
rect 401782 527031 401838 527040
rect 401796 526454 401824 527031
rect 401784 526448 401836 526454
rect 401784 526390 401836 526396
rect 401600 521008 401652 521014
rect 401598 520976 401600 520985
rect 401652 520976 401654 520985
rect 401598 520911 401654 520920
rect 401600 520192 401652 520198
rect 401598 520160 401600 520169
rect 401652 520160 401654 520169
rect 401598 520095 401654 520104
rect 401600 516112 401652 516118
rect 401598 516080 401600 516089
rect 401652 516080 401654 516089
rect 401598 516015 401654 516024
rect 401598 513904 401654 513913
rect 401598 513839 401654 513848
rect 400864 503736 400916 503742
rect 400864 503678 400916 503684
rect 400772 499384 400824 499390
rect 400772 499326 400824 499332
rect 399300 498160 399352 498166
rect 399300 498102 399352 498108
rect 396724 498092 396776 498098
rect 396724 498034 396776 498040
rect 398840 494828 398892 494834
rect 398840 494770 398892 494776
rect 396172 21480 396224 21486
rect 396172 21422 396224 21428
rect 396080 8288 396132 8294
rect 396080 8230 396132 8236
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396184 354 396212 21422
rect 398852 3194 398880 494770
rect 400876 239426 400904 503678
rect 401612 499186 401640 513839
rect 401692 503668 401744 503674
rect 401692 503610 401744 503616
rect 401704 503305 401732 503610
rect 401690 503296 401746 503305
rect 401690 503231 401746 503240
rect 401796 503146 401824 526390
rect 401888 510513 401916 529926
rect 401968 528352 402020 528358
rect 401968 528294 402020 528300
rect 401980 527785 402008 528294
rect 401966 527776 402022 527785
rect 401966 527711 402022 527720
rect 402072 517449 402100 550530
rect 402058 517440 402114 517449
rect 402058 517375 402114 517384
rect 401966 515536 402022 515545
rect 401966 515471 402022 515480
rect 401874 510504 401930 510513
rect 401874 510439 401930 510448
rect 401874 508464 401930 508473
rect 401874 508399 401930 508408
rect 401704 503118 401824 503146
rect 401704 499254 401732 503118
rect 401888 503010 401916 508399
rect 401796 502982 401916 503010
rect 401796 499361 401824 502982
rect 401874 500304 401930 500313
rect 401874 500239 401930 500248
rect 401888 499594 401916 500239
rect 401876 499588 401928 499594
rect 401876 499530 401928 499536
rect 401782 499352 401838 499361
rect 401782 499287 401838 499296
rect 401692 499248 401744 499254
rect 401692 499190 401744 499196
rect 401600 499180 401652 499186
rect 401600 499122 401652 499128
rect 401980 499118 402008 515471
rect 402058 513496 402114 513505
rect 402058 513431 402114 513440
rect 402072 500886 402100 513431
rect 402164 506025 402192 561070
rect 402244 526788 402296 526794
rect 402244 526730 402296 526736
rect 402256 526425 402284 526730
rect 402242 526416 402298 526425
rect 402242 526351 402298 526360
rect 402244 525360 402296 525366
rect 402244 525302 402296 525308
rect 402256 525065 402284 525302
rect 402242 525056 402298 525065
rect 402242 524991 402298 525000
rect 402348 512009 402376 639202
rect 402520 639056 402572 639062
rect 402520 638998 402572 639004
rect 402428 549908 402480 549914
rect 402428 549850 402480 549856
rect 402440 532545 402468 549850
rect 402426 532536 402482 532545
rect 402426 532471 402482 532480
rect 402428 525768 402480 525774
rect 402428 525710 402480 525716
rect 402440 512825 402468 525710
rect 402532 518265 402560 638998
rect 403072 554804 403124 554810
rect 403072 554746 403124 554752
rect 402980 551472 403032 551478
rect 402980 551414 403032 551420
rect 402992 538214 403020 551414
rect 403084 546417 403112 554746
rect 403070 546408 403126 546417
rect 403070 546343 403126 546352
rect 402992 538186 403112 538214
rect 403084 534074 403112 538186
rect 402992 534046 403112 534074
rect 402886 530360 402942 530369
rect 402886 530295 402942 530304
rect 402900 530058 402928 530295
rect 402888 530052 402940 530058
rect 402888 529994 402940 530000
rect 402886 529000 402942 529009
rect 402886 528935 402942 528944
rect 402900 528630 402928 528935
rect 402888 528624 402940 528630
rect 402888 528566 402940 528572
rect 402886 528456 402942 528465
rect 402992 528442 403020 534046
rect 403176 528873 403204 642466
rect 403624 634840 403676 634846
rect 403624 634782 403676 634788
rect 403636 600302 403664 634782
rect 403624 600296 403676 600302
rect 403624 600238 403676 600244
rect 403256 598324 403308 598330
rect 403256 598266 403308 598272
rect 403162 528864 403218 528873
rect 403162 528799 403218 528808
rect 402942 528414 403020 528442
rect 402886 528391 402942 528400
rect 403268 524414 403296 598266
rect 403348 598256 403400 598262
rect 403348 598198 403400 598204
rect 403360 536246 403388 598198
rect 403440 551336 403492 551342
rect 403440 551278 403492 551284
rect 403348 536240 403400 536246
rect 403348 536182 403400 536188
rect 402900 524386 403296 524414
rect 402900 524113 402928 524386
rect 402886 524104 402942 524113
rect 402886 524039 402942 524048
rect 402886 521792 402942 521801
rect 402886 521727 402942 521736
rect 402900 521694 402928 521727
rect 402888 521688 402940 521694
rect 402888 521630 402940 521636
rect 402518 518256 402574 518265
rect 402518 518191 402574 518200
rect 402610 516216 402666 516225
rect 402610 516151 402612 516160
rect 402664 516151 402666 516160
rect 402612 516122 402664 516128
rect 403452 516118 403480 551278
rect 403532 551064 403584 551070
rect 403532 551006 403584 551012
rect 403544 521014 403572 551006
rect 403532 521008 403584 521014
rect 403532 520950 403584 520956
rect 403440 516112 403492 516118
rect 403440 516054 403492 516060
rect 402520 513256 402572 513262
rect 402518 513224 402520 513233
rect 402572 513224 402574 513233
rect 402518 513159 402574 513168
rect 402426 512816 402482 512825
rect 402426 512751 402482 512760
rect 402334 512000 402390 512009
rect 402334 511935 402390 511944
rect 402886 510776 402942 510785
rect 402886 510711 402942 510720
rect 402900 510678 402928 510711
rect 402888 510672 402940 510678
rect 402888 510614 402940 510620
rect 402886 509552 402942 509561
rect 402886 509487 402942 509496
rect 402900 509386 402928 509487
rect 402888 509380 402940 509386
rect 402888 509322 402940 509328
rect 402244 506456 402296 506462
rect 402242 506424 402244 506433
rect 402296 506424 402298 506433
rect 402242 506359 402298 506368
rect 402150 506016 402206 506025
rect 402150 505951 402206 505960
rect 402244 501016 402296 501022
rect 402244 500958 402296 500964
rect 402060 500880 402112 500886
rect 402060 500822 402112 500828
rect 401968 499112 402020 499118
rect 401968 499054 402020 499060
rect 400864 239420 400916 239426
rect 400864 239362 400916 239368
rect 402256 18630 402284 500958
rect 403728 499526 403756 670686
rect 405096 662584 405148 662590
rect 405096 662526 405148 662532
rect 403808 662448 403860 662454
rect 403808 662390 403860 662396
rect 403820 520198 403848 662390
rect 405004 641776 405056 641782
rect 405004 641718 405056 641724
rect 403900 638988 403952 638994
rect 403900 638930 403952 638936
rect 403808 520192 403860 520198
rect 403808 520134 403860 520140
rect 403716 499520 403768 499526
rect 403716 499462 403768 499468
rect 403912 498166 403940 638930
rect 404728 599208 404780 599214
rect 404728 599150 404780 599156
rect 404636 598392 404688 598398
rect 404636 598334 404688 598340
rect 404360 557592 404412 557598
rect 404360 557534 404412 557540
rect 404372 533798 404400 557534
rect 404452 551404 404504 551410
rect 404452 551346 404504 551352
rect 404360 533792 404412 533798
rect 404360 533734 404412 533740
rect 404464 531282 404492 551346
rect 404544 550860 404596 550866
rect 404544 550802 404596 550808
rect 404556 543454 404584 550802
rect 404544 543448 404596 543454
rect 404544 543390 404596 543396
rect 404452 531276 404504 531282
rect 404452 531218 404504 531224
rect 404648 528358 404676 598334
rect 404740 531962 404768 599150
rect 405016 599146 405044 641718
rect 405004 599140 405056 599146
rect 405004 599082 405056 599088
rect 404820 554056 404872 554062
rect 404820 553998 404872 554004
rect 404728 531956 404780 531962
rect 404728 531898 404780 531904
rect 404636 528352 404688 528358
rect 404636 528294 404688 528300
rect 404832 506462 404860 553998
rect 404912 550724 404964 550730
rect 404912 550666 404964 550672
rect 404924 525366 404952 550666
rect 405108 526794 405136 662526
rect 405740 662516 405792 662522
rect 405740 662458 405792 662464
rect 405280 642184 405332 642190
rect 405280 642126 405332 642132
rect 405188 642048 405240 642054
rect 405188 641990 405240 641996
rect 405096 526788 405148 526794
rect 405096 526730 405148 526736
rect 405096 525836 405148 525842
rect 405096 525778 405148 525784
rect 404912 525360 404964 525366
rect 404912 525302 404964 525308
rect 404910 509416 404966 509425
rect 404910 509351 404912 509360
rect 404964 509351 404966 509360
rect 404912 509322 404964 509328
rect 404820 506456 404872 506462
rect 404820 506398 404872 506404
rect 405004 505164 405056 505170
rect 405004 505106 405056 505112
rect 403900 498160 403952 498166
rect 403900 498102 403952 498108
rect 402980 493400 403032 493406
rect 402980 493342 403032 493348
rect 402244 18624 402296 18630
rect 402244 18566 402296 18572
rect 402992 16574 403020 493342
rect 405016 18698 405044 505106
rect 405108 280090 405136 525778
rect 405200 498098 405228 641990
rect 405188 498092 405240 498098
rect 405188 498034 405240 498040
rect 405292 498030 405320 642126
rect 405752 513262 405780 662458
rect 405832 661360 405884 661366
rect 405832 661302 405884 661308
rect 405740 513256 405792 513262
rect 405740 513198 405792 513204
rect 405844 503674 405872 661302
rect 406396 529922 406424 700266
rect 407120 530528 407172 530534
rect 407120 530470 407172 530476
rect 406384 529916 406436 529922
rect 406384 529858 406436 529864
rect 405924 516180 405976 516186
rect 405924 516122 405976 516128
rect 405832 503668 405884 503674
rect 405832 503610 405884 503616
rect 405280 498024 405332 498030
rect 405280 497966 405332 497972
rect 405096 280084 405148 280090
rect 405096 280026 405148 280032
rect 405004 18692 405056 18698
rect 405004 18634 405056 18640
rect 405936 16574 405964 516122
rect 407132 16574 407160 530470
rect 409880 530120 409932 530126
rect 409880 530062 409932 530068
rect 409144 528624 409196 528630
rect 409144 528566 409196 528572
rect 409156 167006 409184 528566
rect 409144 167000 409196 167006
rect 409144 166942 409196 166948
rect 408500 89072 408552 89078
rect 408500 89014 408552 89020
rect 408512 16574 408540 89014
rect 409892 16574 409920 530062
rect 412652 513330 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 422944 661836 422996 661842
rect 422944 661778 422996 661784
rect 418804 552288 418856 552294
rect 418804 552230 418856 552236
rect 414664 552152 414716 552158
rect 414664 552094 414716 552100
rect 412640 513324 412692 513330
rect 412640 513266 412692 513272
rect 414020 497548 414072 497554
rect 414020 497490 414072 497496
rect 412640 491972 412692 491978
rect 412640 491914 412692 491920
rect 402992 16546 403664 16574
rect 405936 16546 406056 16574
rect 407132 16546 407252 16574
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 402520 8288 402572 8294
rect 402520 8230 402572 8236
rect 398840 3188 398892 3194
rect 398840 3130 398892 3136
rect 400128 3188 400180 3194
rect 400128 3130 400180 3136
rect 400140 480 400168 3130
rect 402532 480 402560 8230
rect 403636 480 403664 16546
rect 406028 480 406056 16546
rect 407224 480 407252 16546
rect 396510 354 396622 480
rect 396184 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 491914
rect 414032 16574 414060 497490
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 414676 3398 414704 552094
rect 416780 531888 416832 531894
rect 416780 531830 416832 531836
rect 416044 528624 416096 528630
rect 416044 528566 416096 528572
rect 415400 89004 415452 89010
rect 415400 88946 415452 88952
rect 414664 3392 414716 3398
rect 414664 3334 414716 3340
rect 415412 3194 415440 88946
rect 416056 35222 416084 528566
rect 416044 35216 416096 35222
rect 416044 35158 416096 35164
rect 416792 16574 416820 531830
rect 418816 206990 418844 552230
rect 420184 552084 420236 552090
rect 420184 552026 420236 552032
rect 418804 206984 418856 206990
rect 418804 206926 418856 206932
rect 418804 63572 418856 63578
rect 418804 63514 418856 63520
rect 416792 16546 417464 16574
rect 415400 3188 415452 3194
rect 415400 3130 415452 3136
rect 416688 3188 416740 3194
rect 416688 3130 416740 3136
rect 416700 480 416728 3130
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 418816 7818 418844 63514
rect 420196 17338 420224 552026
rect 420920 527196 420972 527202
rect 420920 527138 420972 527144
rect 420184 17332 420236 17338
rect 420184 17274 420236 17280
rect 418804 7812 418856 7818
rect 418804 7754 418856 7760
rect 420184 3392 420236 3398
rect 420184 3334 420236 3340
rect 420196 480 420224 3334
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 527138
rect 422956 525774 422984 661778
rect 430580 552220 430632 552226
rect 430580 552162 430632 552168
rect 422944 525768 422996 525774
rect 422944 525710 422996 525716
rect 423680 521688 423732 521694
rect 423680 521630 423732 521636
rect 422944 509312 422996 509318
rect 422944 509254 422996 509260
rect 422956 21486 422984 509254
rect 422944 21480 422996 21486
rect 422944 21422 422996 21428
rect 423692 3210 423720 521630
rect 427820 497684 427872 497690
rect 427820 497626 427872 497632
rect 426440 177336 426492 177342
rect 426440 177278 426492 177284
rect 423772 21480 423824 21486
rect 423772 21422 423824 21428
rect 423784 3398 423812 21422
rect 426452 16574 426480 177278
rect 427832 16574 427860 497626
rect 430592 16574 430620 552162
rect 444380 551540 444432 551546
rect 444380 551482 444432 551488
rect 437480 541000 437532 541006
rect 437480 540942 437532 540948
rect 434720 531956 434772 531962
rect 434720 531898 434772 531904
rect 433340 499588 433392 499594
rect 433340 499530 433392 499536
rect 431960 352572 432012 352578
rect 431960 352514 432012 352520
rect 431972 16574 432000 352514
rect 433352 16574 433380 499530
rect 434732 16574 434760 531898
rect 436744 517540 436796 517546
rect 436744 517482 436796 517488
rect 436756 36582 436784 517482
rect 436836 503804 436888 503810
rect 436836 503746 436888 503752
rect 436848 224330 436876 503746
rect 436836 224324 436888 224330
rect 436836 224266 436888 224272
rect 436744 36576 436796 36582
rect 436744 36518 436796 36524
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 431972 16546 432092 16574
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 423772 3392 423824 3398
rect 423772 3334 423824 3340
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 423692 3182 423812 3210
rect 423784 480 423812 3182
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 430868 480 430896 16546
rect 432064 480 432092 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 540942
rect 438860 531820 438912 531826
rect 438860 531762 438912 531768
rect 438872 16574 438900 531762
rect 441620 513392 441672 513398
rect 441620 513334 441672 513340
rect 440884 502376 440936 502382
rect 440884 502318 440936 502324
rect 440896 22778 440924 502318
rect 440884 22772 440936 22778
rect 440884 22714 440936 22720
rect 441632 16574 441660 513334
rect 438872 16546 439176 16574
rect 441632 16546 442672 16574
rect 439148 480 439176 16546
rect 440240 15972 440292 15978
rect 440240 15914 440292 15920
rect 440252 3194 440280 15914
rect 440240 3188 440292 3194
rect 440240 3130 440292 3136
rect 441528 3188 441580 3194
rect 441528 3130 441580 3136
rect 441540 480 441568 3130
rect 442644 480 442672 16546
rect 444392 6914 444420 551482
rect 448520 531548 448572 531554
rect 448520 531490 448572 531496
rect 445024 509380 445076 509386
rect 445024 509322 445076 509328
rect 445036 9110 445064 509322
rect 445760 494896 445812 494902
rect 445760 494838 445812 494844
rect 445024 9104 445076 9110
rect 445024 9046 445076 9052
rect 444392 6886 445064 6914
rect 445036 480 445064 6886
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 494838
rect 448532 3398 448560 531490
rect 458180 530052 458232 530058
rect 458180 529994 458232 530000
rect 456800 523048 456852 523054
rect 456800 522990 456852 522996
rect 450544 520328 450596 520334
rect 450544 520270 450596 520276
rect 448610 177304 448666 177313
rect 448610 177239 448666 177248
rect 448520 3392 448572 3398
rect 448520 3334 448572 3340
rect 448624 480 448652 177239
rect 450556 18766 450584 520270
rect 454684 518968 454736 518974
rect 454684 518910 454736 518916
rect 451280 510672 451332 510678
rect 451280 510614 451332 510620
rect 450544 18760 450596 18766
rect 450544 18702 450596 18708
rect 451292 16574 451320 510614
rect 454696 17270 454724 518910
rect 454684 17264 454736 17270
rect 454684 17206 454736 17212
rect 456812 16574 456840 522990
rect 458192 16574 458220 529994
rect 460204 513460 460256 513466
rect 460204 513402 460256 513408
rect 459560 497616 459612 497622
rect 459560 497558 459612 497564
rect 459572 16574 459600 497558
rect 460216 478174 460244 513402
rect 462332 510610 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477040 700528 477092 700534
rect 477040 700470 477092 700476
rect 475752 665848 475804 665854
rect 475752 665790 475804 665796
rect 475660 661700 475712 661706
rect 475660 661642 475712 661648
rect 472624 641844 472676 641850
rect 472624 641786 472676 641792
rect 472636 599078 472664 641786
rect 472624 599072 472676 599078
rect 472624 599014 472676 599020
rect 471244 598256 471296 598262
rect 471244 598198 471296 598204
rect 463700 531616 463752 531622
rect 463700 531558 463752 531564
rect 462964 510672 463016 510678
rect 462964 510614 463016 510620
rect 462320 510604 462372 510610
rect 462320 510546 462372 510552
rect 460204 478168 460256 478174
rect 460204 478110 460256 478116
rect 462976 37942 463004 510614
rect 462964 37936 463016 37942
rect 462964 37878 463016 37884
rect 463712 16574 463740 531558
rect 468484 530324 468536 530330
rect 468484 530266 468536 530272
rect 466460 517608 466512 517614
rect 466460 517550 466512 517556
rect 466472 16574 466500 517550
rect 451292 16546 451688 16574
rect 456812 16546 456932 16574
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 463712 16546 464016 16574
rect 466472 16546 467512 16574
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 449820 480 449848 3334
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 455696 11756 455748 11762
rect 455696 11698 455748 11704
rect 453304 3664 453356 3670
rect 453304 3606 453356 3612
rect 453316 480 453344 3606
rect 455708 480 455736 11698
rect 456904 480 456932 16546
rect 459204 480 459232 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 463988 480 464016 16546
rect 467484 480 467512 16546
rect 468496 3466 468524 530266
rect 468576 499588 468628 499594
rect 468576 499530 468628 499536
rect 468588 250510 468616 499530
rect 471256 499458 471284 598198
rect 474002 579048 474058 579057
rect 474002 578983 474058 578992
rect 473360 531412 473412 531418
rect 473360 531354 473412 531360
rect 472624 530256 472676 530262
rect 472624 530198 472676 530204
rect 471336 523252 471388 523258
rect 471336 523194 471388 523200
rect 471244 499452 471296 499458
rect 471244 499394 471296 499400
rect 470600 497820 470652 497826
rect 470600 497762 470652 497768
rect 468576 250504 468628 250510
rect 468576 250446 468628 250452
rect 468484 3460 468536 3466
rect 468484 3402 468536 3408
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 497762
rect 471348 479534 471376 523194
rect 471336 479528 471388 479534
rect 471336 479470 471388 479476
rect 472636 3534 472664 530198
rect 472716 505572 472768 505578
rect 472716 505514 472768 505520
rect 472728 45558 472756 505514
rect 472716 45552 472768 45558
rect 472716 45494 472768 45500
rect 473372 16574 473400 531354
rect 474016 498098 474044 578983
rect 475476 532024 475528 532030
rect 475476 531966 475528 531972
rect 475384 531752 475436 531758
rect 475384 531694 475436 531700
rect 474004 498092 474056 498098
rect 474004 498034 474056 498040
rect 473372 16546 474136 16574
rect 473452 5024 473504 5030
rect 473452 4966 473504 4972
rect 472624 3528 472676 3534
rect 472624 3470 472676 3476
rect 473464 480 473492 4966
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475396 7750 475424 531694
rect 475488 21418 475516 531966
rect 475568 530460 475620 530466
rect 475568 530402 475620 530408
rect 475580 117298 475608 530402
rect 475672 498166 475700 661642
rect 475764 525638 475792 665790
rect 475844 550656 475896 550662
rect 475844 550598 475896 550604
rect 475752 525632 475804 525638
rect 475752 525574 475804 525580
rect 475660 498160 475712 498166
rect 475660 498102 475712 498108
rect 475856 498030 475884 550598
rect 476764 531684 476816 531690
rect 476764 531626 476816 531632
rect 475844 498024 475896 498030
rect 475844 497966 475896 497972
rect 475568 117292 475620 117298
rect 475568 117234 475620 117240
rect 475476 21412 475528 21418
rect 475476 21354 475528 21360
rect 476776 13122 476804 531626
rect 476948 531480 477000 531486
rect 476948 531422 477000 531428
rect 476856 531344 476908 531350
rect 476856 531286 476908 531292
rect 476868 31074 476896 531286
rect 476960 225622 476988 531422
rect 477052 499390 477080 700470
rect 477132 698964 477184 698970
rect 477132 698906 477184 698912
rect 477144 517478 477172 698906
rect 477224 659864 477276 659870
rect 477224 659806 477276 659812
rect 477132 517472 477184 517478
rect 477132 517414 477184 517420
rect 477040 499384 477092 499390
rect 477040 499326 477092 499332
rect 477236 497962 477264 659806
rect 477512 654134 477540 702406
rect 527192 699718 527220 703520
rect 543476 700398 543504 703520
rect 559668 700466 559696 703520
rect 559656 700460 559708 700466
rect 559656 700402 559708 700408
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 520924 699712 520976 699718
rect 520924 699654 520976 699660
rect 527180 699712 527232 699718
rect 527180 699654 527232 699660
rect 512000 661292 512052 661298
rect 512000 661234 512052 661240
rect 478880 661224 478932 661230
rect 512012 661201 512040 661234
rect 478880 661166 478932 661172
rect 511998 661192 512054 661201
rect 477512 654106 477632 654134
rect 477604 625154 477632 654106
rect 478694 636168 478750 636177
rect 478694 636103 478750 636112
rect 478708 634846 478736 636103
rect 478696 634840 478748 634846
rect 478696 634782 478748 634788
rect 477512 625126 477632 625154
rect 477512 536110 477540 625126
rect 478142 617808 478198 617817
rect 478142 617743 478198 617752
rect 478156 598806 478184 617743
rect 478144 598800 478196 598806
rect 478144 598742 478196 598748
rect 478892 538214 478920 661166
rect 484400 661156 484452 661162
rect 511998 661127 512054 661136
rect 484400 661098 484452 661104
rect 484412 661065 484440 661098
rect 498200 661088 498252 661094
rect 484398 661056 484454 661065
rect 484398 660991 484454 661000
rect 498198 661056 498200 661065
rect 498252 661056 498254 661065
rect 498198 660991 498254 661000
rect 488540 660476 488592 660482
rect 488540 660418 488592 660424
rect 488552 660249 488580 660418
rect 500960 660340 501012 660346
rect 500960 660282 501012 660288
rect 488538 660240 488594 660249
rect 488538 660175 488594 660184
rect 500972 659841 501000 660282
rect 500958 659832 501014 659841
rect 500958 659767 501014 659776
rect 493232 641844 493284 641850
rect 493232 641786 493284 641792
rect 493244 639962 493272 641786
rect 510620 641776 510672 641782
rect 510620 641718 510672 641724
rect 510632 639962 510660 641718
rect 493244 639934 493580 639962
rect 510632 639934 510968 639962
rect 479720 600086 480056 600114
rect 496464 600086 496800 600114
rect 513852 600086 514188 600114
rect 479720 596873 479748 600086
rect 496464 598262 496492 600086
rect 513852 598874 513880 600086
rect 513840 598868 513892 598874
rect 513840 598810 513892 598816
rect 496452 598256 496504 598262
rect 496452 598198 496504 598204
rect 479706 596864 479762 596873
rect 479706 596799 479762 596808
rect 510712 595468 510764 595474
rect 510712 595410 510764 595416
rect 499580 594108 499632 594114
rect 499580 594050 499632 594056
rect 498200 592680 498252 592686
rect 498200 592622 498252 592628
rect 485872 590708 485924 590714
rect 485872 590650 485924 590656
rect 483112 559564 483164 559570
rect 483112 559506 483164 559512
rect 478892 538186 479656 538214
rect 477500 536104 477552 536110
rect 477500 536046 477552 536052
rect 478880 530392 478932 530398
rect 478880 530334 478932 530340
rect 477500 529916 477552 529922
rect 477500 529858 477552 529864
rect 477512 529689 477540 529858
rect 477498 529680 477554 529689
rect 477498 529615 477554 529624
rect 477500 528624 477552 528630
rect 477498 528592 477500 528601
rect 477552 528592 477554 528601
rect 477498 528527 477554 528536
rect 477498 527232 477554 527241
rect 477498 527167 477500 527176
rect 477552 527167 477554 527176
rect 477500 527138 477552 527144
rect 478892 526454 478920 530334
rect 479628 529938 479656 538186
rect 481548 533384 481600 533390
rect 481548 533326 481600 533332
rect 480996 530052 481048 530058
rect 480996 529994 481048 530000
rect 481008 529938 481036 529994
rect 481560 529938 481588 533326
rect 481822 532672 481878 532681
rect 481822 532607 481878 532616
rect 479628 529910 480056 529938
rect 480700 529910 481036 529938
rect 481344 529910 481588 529938
rect 481836 529938 481864 532607
rect 482926 529952 482982 529961
rect 481836 529910 481988 529938
rect 482632 529910 482926 529938
rect 483124 529938 483152 559506
rect 485884 538214 485912 590650
rect 498212 538214 498240 592622
rect 485884 538186 486096 538214
rect 498212 538186 498332 538214
rect 485504 536852 485556 536858
rect 485504 536794 485556 536800
rect 484674 532672 484730 532681
rect 484674 532607 484730 532616
rect 483572 531344 483624 531350
rect 483572 531286 483624 531292
rect 483584 529938 483612 531286
rect 484688 529938 484716 532607
rect 485044 530596 485096 530602
rect 485044 530538 485096 530544
rect 485056 530330 485084 530538
rect 485044 530324 485096 530330
rect 485044 530266 485096 530272
rect 485516 529938 485544 536794
rect 485826 530188 485878 530194
rect 485826 530130 485878 530136
rect 483124 529910 483276 529938
rect 483584 529910 483920 529938
rect 484564 529910 484716 529938
rect 485208 529910 485544 529938
rect 485838 529924 485866 530130
rect 486068 529938 486096 538186
rect 488998 532672 489054 532681
rect 488998 532607 489054 532616
rect 487436 531548 487488 531554
rect 487436 531490 487488 531496
rect 486792 531412 486844 531418
rect 486792 531354 486844 531360
rect 486804 529938 486832 531354
rect 487448 529938 487476 531490
rect 488080 531480 488132 531486
rect 488080 531422 488132 531428
rect 488092 529938 488120 531422
rect 489012 529938 489040 532607
rect 492680 532024 492732 532030
rect 492680 531966 492732 531972
rect 494428 532024 494480 532030
rect 494428 531966 494480 531972
rect 491944 530596 491996 530602
rect 491944 530538 491996 530544
rect 491622 530120 491674 530126
rect 491622 530062 491674 530068
rect 491208 529984 491260 529990
rect 486068 529910 486496 529938
rect 486804 529910 487140 529938
rect 487448 529910 487784 529938
rect 488092 529910 488428 529938
rect 489012 529910 489072 529938
rect 491004 529932 491208 529938
rect 491004 529926 491260 529932
rect 491004 529910 491248 529926
rect 491634 529924 491662 530062
rect 491956 529938 491984 530538
rect 492692 529938 492720 531966
rect 493876 531412 493928 531418
rect 493876 531354 493928 531360
rect 493888 529938 493916 531354
rect 494440 529938 494468 531966
rect 497740 531888 497792 531894
rect 497740 531830 497792 531836
rect 496452 531820 496504 531826
rect 496452 531762 496504 531768
rect 495440 531616 495492 531622
rect 495440 531558 495492 531564
rect 494520 530460 494572 530466
rect 494520 530402 494572 530408
rect 491956 529910 492292 529938
rect 492692 529910 492936 529938
rect 493580 529910 493916 529938
rect 494224 529910 494468 529938
rect 494532 529938 494560 530402
rect 495452 529938 495480 531558
rect 495808 530528 495860 530534
rect 495808 530470 495860 530476
rect 495820 529938 495848 530470
rect 496464 529938 496492 531762
rect 497096 530256 497148 530262
rect 497096 530198 497148 530204
rect 497108 529938 497136 530198
rect 497752 529938 497780 531830
rect 498304 529938 498332 538186
rect 499304 531616 499356 531622
rect 499304 531558 499356 531564
rect 499316 529938 499344 531558
rect 499592 529938 499620 594050
rect 506480 585812 506532 585818
rect 506480 585754 506532 585760
rect 506492 538214 506520 585754
rect 506492 538186 507348 538214
rect 502892 536104 502944 536110
rect 502892 536046 502944 536052
rect 501878 532672 501934 532681
rect 501878 532607 501934 532616
rect 500958 532536 501014 532545
rect 500958 532471 501014 532480
rect 500316 530392 500368 530398
rect 500316 530334 500368 530340
rect 500328 529938 500356 530334
rect 500972 529938 501000 532471
rect 501892 529938 501920 532607
rect 502904 529938 502932 536046
rect 505560 531956 505612 531962
rect 505560 531898 505612 531904
rect 504180 531548 504232 531554
rect 504180 531490 504232 531496
rect 504192 529938 504220 531490
rect 505468 531344 505520 531350
rect 505468 531286 505520 531292
rect 505480 529938 505508 531286
rect 494532 529910 494868 529938
rect 495452 529910 495512 529938
rect 495820 529910 496156 529938
rect 496464 529910 496800 529938
rect 497108 529910 497444 529938
rect 497752 529910 498088 529938
rect 498304 529910 498732 529938
rect 499316 529910 499376 529938
rect 499592 529910 500020 529938
rect 500328 529910 500664 529938
rect 500972 529910 501308 529938
rect 501892 529910 501952 529938
rect 502904 529910 503240 529938
rect 503884 529910 504220 529938
rect 505172 529910 505508 529938
rect 505572 529938 505600 531898
rect 506112 531752 506164 531758
rect 506112 531694 506164 531700
rect 507216 531752 507268 531758
rect 507216 531694 507268 531700
rect 506124 529938 506152 531694
rect 507228 529938 507256 531694
rect 505572 529910 505816 529938
rect 506124 529910 506460 529938
rect 507104 529910 507256 529938
rect 507320 529938 507348 538186
rect 508780 531684 508832 531690
rect 508780 531626 508832 531632
rect 508688 531480 508740 531486
rect 508688 531422 508740 531428
rect 508700 529938 508728 531422
rect 507320 529910 507748 529938
rect 508392 529910 508728 529938
rect 508792 529938 508820 531626
rect 509884 531412 509936 531418
rect 509884 531354 509936 531360
rect 508792 529910 509036 529938
rect 482926 529887 482982 529896
rect 489550 529544 489606 529553
rect 502430 529544 502486 529553
rect 489606 529502 489716 529530
rect 489550 529479 489606 529488
rect 504178 529544 504234 529553
rect 502486 529502 502596 529530
rect 502430 529479 502486 529488
rect 504234 529502 504528 529530
rect 504178 529479 504234 529488
rect 509680 529230 509832 529258
rect 509804 528902 509832 529230
rect 509792 528896 509844 528902
rect 509792 528838 509844 528844
rect 509896 527882 509924 531354
rect 510620 531344 510672 531350
rect 510620 531286 510672 531292
rect 509884 527876 509936 527882
rect 509884 527818 509936 527824
rect 479154 527504 479210 527513
rect 479154 527439 479210 527448
rect 478880 526448 478932 526454
rect 478880 526390 478932 526396
rect 479062 526144 479118 526153
rect 479062 526079 479118 526088
rect 477498 525872 477554 525881
rect 477498 525807 477500 525816
rect 477552 525807 477554 525816
rect 477500 525778 477552 525784
rect 478696 525768 478748 525774
rect 478696 525710 478748 525716
rect 477960 525632 478012 525638
rect 477958 525600 477960 525609
rect 478012 525600 478014 525609
rect 477958 525535 478014 525544
rect 478708 525065 478736 525710
rect 478694 525056 478750 525065
rect 478694 524991 478750 525000
rect 477498 523424 477554 523433
rect 477498 523359 477554 523368
rect 477512 523258 477540 523359
rect 477500 523252 477552 523258
rect 477500 523194 477552 523200
rect 477498 523152 477554 523161
rect 477498 523087 477554 523096
rect 477512 523054 477540 523087
rect 477500 523048 477552 523054
rect 477500 522990 477552 522996
rect 478418 522064 478474 522073
rect 478418 521999 478474 522008
rect 477958 521792 478014 521801
rect 477958 521727 478014 521736
rect 477498 520704 477554 520713
rect 477498 520639 477554 520648
rect 477512 520334 477540 520639
rect 477500 520328 477552 520334
rect 477500 520270 477552 520276
rect 477590 517984 477646 517993
rect 477590 517919 477646 517928
rect 477498 517712 477554 517721
rect 477498 517647 477554 517656
rect 477512 517546 477540 517647
rect 477604 517614 477632 517919
rect 477592 517608 477644 517614
rect 477592 517550 477644 517556
rect 477500 517540 477552 517546
rect 477500 517482 477552 517488
rect 477590 513904 477646 513913
rect 477590 513839 477646 513848
rect 477498 513496 477554 513505
rect 477604 513466 477632 513839
rect 477498 513431 477554 513440
rect 477592 513460 477644 513466
rect 477512 513398 477540 513431
rect 477592 513402 477644 513408
rect 477500 513392 477552 513398
rect 477500 513334 477552 513340
rect 477592 513324 477644 513330
rect 477592 513266 477644 513272
rect 477604 512825 477632 513266
rect 477590 512816 477646 512825
rect 477590 512751 477646 512760
rect 477590 511184 477646 511193
rect 477590 511119 477646 511128
rect 477604 510678 477632 511119
rect 477592 510672 477644 510678
rect 477592 510614 477644 510620
rect 477866 510640 477922 510649
rect 477500 510604 477552 510610
rect 477866 510575 477922 510584
rect 477500 510546 477552 510552
rect 477512 510513 477540 510546
rect 477498 510504 477554 510513
rect 477498 510439 477554 510448
rect 477498 509416 477554 509425
rect 477498 509351 477554 509360
rect 477512 509318 477540 509351
rect 477500 509312 477552 509318
rect 477500 509254 477552 509260
rect 477498 505744 477554 505753
rect 477498 505679 477554 505688
rect 477512 505578 477540 505679
rect 477500 505572 477552 505578
rect 477500 505514 477552 505520
rect 477498 505336 477554 505345
rect 477498 505271 477554 505280
rect 477512 505170 477540 505271
rect 477500 505164 477552 505170
rect 477500 505106 477552 505112
rect 477590 504384 477646 504393
rect 477590 504319 477646 504328
rect 477498 503976 477554 503985
rect 477498 503911 477554 503920
rect 477512 503742 477540 503911
rect 477604 503810 477632 504319
rect 477592 503804 477644 503810
rect 477592 503746 477644 503752
rect 477500 503736 477552 503742
rect 477500 503678 477552 503684
rect 477498 502616 477554 502625
rect 477498 502551 477554 502560
rect 477512 502382 477540 502551
rect 477500 502376 477552 502382
rect 477500 502318 477552 502324
rect 477498 501664 477554 501673
rect 477498 501599 477554 501608
rect 477512 501022 477540 501599
rect 477500 501016 477552 501022
rect 477500 500958 477552 500964
rect 477498 500168 477554 500177
rect 477498 500103 477554 500112
rect 477512 499594 477540 500103
rect 477500 499588 477552 499594
rect 477500 499530 477552 499536
rect 477224 497956 477276 497962
rect 477224 497898 477276 497904
rect 476948 225616 477000 225622
rect 476948 225558 477000 225564
rect 477880 177410 477908 510575
rect 477868 177404 477920 177410
rect 477868 177346 477920 177352
rect 476856 31068 476908 31074
rect 476856 31010 476908 31016
rect 476764 13116 476816 13122
rect 476764 13058 476816 13064
rect 477868 10328 477920 10334
rect 477868 10270 477920 10276
rect 475384 7744 475436 7750
rect 475384 7686 475436 7692
rect 477880 3482 477908 10270
rect 477972 5030 478000 521727
rect 478234 517032 478290 517041
rect 478234 516967 478290 516976
rect 478142 507104 478198 507113
rect 478142 507039 478198 507048
rect 478156 280158 478184 507039
rect 478248 496806 478276 516967
rect 478432 502806 478460 521999
rect 478602 520296 478658 520305
rect 478602 520231 478658 520240
rect 478510 519344 478566 519353
rect 478510 519279 478566 519288
rect 478524 518974 478552 519279
rect 478512 518968 478564 518974
rect 478512 518910 478564 518916
rect 478512 517472 478564 517478
rect 478512 517414 478564 517420
rect 478524 516905 478552 517414
rect 478510 516896 478566 516905
rect 478510 516831 478566 516840
rect 478510 507920 478566 507929
rect 478510 507855 478566 507864
rect 478340 502778 478460 502806
rect 478236 496800 478288 496806
rect 478236 496742 478288 496748
rect 478340 495446 478368 502778
rect 478524 502738 478552 507855
rect 478432 502710 478552 502738
rect 478432 498234 478460 502710
rect 478512 502648 478564 502654
rect 478512 502590 478564 502596
rect 478420 498228 478472 498234
rect 478420 498170 478472 498176
rect 478328 495440 478380 495446
rect 478328 495382 478380 495388
rect 478144 280152 478196 280158
rect 478144 280094 478196 280100
rect 478524 177342 478552 502590
rect 478616 500954 478644 520231
rect 478694 519072 478750 519081
rect 478694 519007 478750 519016
rect 478604 500948 478656 500954
rect 478604 500890 478656 500896
rect 478512 177336 478564 177342
rect 478512 177278 478564 177284
rect 478708 7750 478736 519007
rect 478970 515264 479026 515273
rect 478970 515199 479026 515208
rect 478786 512952 478842 512961
rect 478786 512887 478842 512896
rect 478800 508502 478828 512887
rect 478788 508496 478840 508502
rect 478788 508438 478840 508444
rect 478786 508328 478842 508337
rect 478786 508263 478842 508272
rect 478800 502654 478828 508263
rect 478788 502648 478840 502654
rect 478788 502590 478840 502596
rect 478786 500984 478842 500993
rect 478786 500919 478842 500928
rect 478800 499526 478828 500919
rect 478788 499520 478840 499526
rect 478788 499462 478840 499468
rect 478984 341562 479012 515199
rect 479076 486470 479104 526079
rect 479168 496262 479196 527439
rect 510632 526561 510660 531286
rect 510618 526552 510674 526561
rect 510618 526487 510674 526496
rect 509882 523016 509938 523025
rect 509882 522951 509938 522960
rect 509790 517984 509846 517993
rect 509790 517919 509846 517928
rect 479246 514856 479302 514865
rect 479246 514791 479302 514800
rect 479260 498778 479288 514791
rect 479524 508496 479576 508502
rect 479524 508438 479576 508444
rect 479430 506560 479486 506569
rect 479430 506495 479486 506504
rect 479338 503024 479394 503033
rect 479338 502959 479394 502968
rect 479248 498772 479300 498778
rect 479248 498714 479300 498720
rect 479156 496256 479208 496262
rect 479156 496198 479208 496204
rect 479352 496126 479380 502959
rect 479340 496120 479392 496126
rect 479340 496062 479392 496068
rect 479064 486464 479116 486470
rect 479064 486406 479116 486412
rect 478972 341556 479024 341562
rect 478972 341498 479024 341504
rect 478696 7744 478748 7750
rect 478696 7686 478748 7692
rect 477960 5024 478012 5030
rect 477960 4966 478012 4972
rect 479444 3534 479472 506495
rect 479536 273222 479564 508438
rect 479720 500126 480056 500154
rect 479720 496194 479748 500126
rect 480686 499882 480714 500140
rect 481330 499882 481358 500140
rect 481974 499882 482002 500140
rect 482618 499882 482646 500140
rect 483262 499882 483290 500140
rect 483906 499882 483934 500140
rect 484550 499882 484578 500140
rect 485194 499882 485222 500140
rect 485838 499882 485866 500140
rect 486482 499882 486510 500140
rect 487126 499882 487154 500140
rect 480640 499854 480714 499882
rect 481284 499854 481358 499882
rect 481928 499854 482002 499882
rect 482572 499854 482646 499882
rect 483216 499854 483290 499882
rect 483860 499854 483934 499882
rect 484504 499854 484578 499882
rect 485148 499854 485222 499882
rect 485792 499854 485866 499882
rect 486436 499854 486510 499882
rect 487080 499854 487154 499882
rect 487770 499882 487798 500140
rect 488414 499882 488442 500140
rect 489058 499882 489086 500140
rect 489702 499882 489730 500140
rect 490346 499882 490374 500140
rect 487770 499854 487844 499882
rect 479708 496188 479760 496194
rect 479708 496130 479760 496136
rect 480640 476814 480668 499854
rect 480904 498228 480956 498234
rect 480904 498170 480956 498176
rect 480628 476808 480680 476814
rect 480628 476750 480680 476756
rect 479524 273216 479576 273222
rect 479524 273158 479576 273164
rect 480352 62144 480404 62150
rect 480352 62086 480404 62092
rect 480364 16574 480392 62086
rect 480916 33114 480944 498170
rect 480996 495440 481048 495446
rect 480996 495382 481048 495388
rect 481008 73166 481036 495382
rect 481088 494012 481140 494018
rect 481088 493954 481140 493960
rect 481100 109002 481128 493954
rect 481088 108996 481140 109002
rect 481088 108938 481140 108944
rect 480996 73160 481048 73166
rect 480996 73102 481048 73108
rect 481284 40798 481312 499854
rect 481640 498772 481692 498778
rect 481640 498714 481692 498720
rect 481272 40792 481324 40798
rect 481272 40734 481324 40740
rect 480904 33108 480956 33114
rect 480904 33050 480956 33056
rect 481652 16574 481680 498714
rect 481928 497418 481956 499854
rect 482376 499520 482428 499526
rect 482376 499462 482428 499468
rect 481916 497412 481968 497418
rect 481916 497354 481968 497360
rect 482284 496800 482336 496806
rect 482284 496742 482336 496748
rect 480364 16546 480576 16574
rect 481652 16546 481772 16574
rect 479432 3528 479484 3534
rect 477880 3454 478184 3482
rect 479432 3470 479484 3476
rect 478156 480 478184 3454
rect 480548 480 480576 16546
rect 481744 480 481772 16546
rect 482296 3466 482324 496742
rect 482388 485790 482416 499462
rect 482376 485784 482428 485790
rect 482376 485726 482428 485732
rect 482572 354006 482600 499854
rect 483216 494766 483244 499854
rect 483204 494760 483256 494766
rect 483204 494702 483256 494708
rect 483860 494018 483888 499854
rect 484504 498166 484532 499854
rect 484492 498160 484544 498166
rect 484492 498102 484544 498108
rect 485148 497826 485176 499854
rect 485136 497820 485188 497826
rect 485136 497762 485188 497768
rect 485044 496868 485096 496874
rect 485044 496810 485096 496816
rect 483848 494012 483900 494018
rect 483848 493954 483900 493960
rect 482560 354000 482612 354006
rect 482560 353942 482612 353948
rect 485056 268462 485084 496810
rect 485792 276690 485820 499854
rect 485780 276684 485832 276690
rect 485780 276626 485832 276632
rect 485044 268456 485096 268462
rect 485044 268398 485096 268404
rect 486436 233238 486464 499854
rect 487080 497486 487108 499854
rect 487816 499458 487844 499854
rect 488368 499854 488442 499882
rect 489012 499854 489086 499882
rect 489656 499854 489730 499882
rect 490300 499854 490374 499882
rect 490990 499882 491018 500140
rect 491634 499882 491662 500140
rect 490990 499854 491064 499882
rect 487804 499452 487856 499458
rect 487804 499394 487856 499400
rect 487068 497480 487120 497486
rect 487068 497422 487120 497428
rect 488368 496874 488396 499854
rect 488356 496868 488408 496874
rect 488356 496810 488408 496816
rect 488632 496256 488684 496262
rect 488632 496198 488684 496204
rect 486424 233232 486476 233238
rect 486424 233174 486476 233180
rect 482376 66292 482428 66298
rect 482376 66234 482428 66240
rect 482388 8294 482416 66234
rect 488644 16574 488672 496198
rect 488644 16546 488856 16574
rect 482376 8288 482428 8294
rect 482376 8230 482428 8236
rect 487620 8288 487672 8294
rect 487620 8230 487672 8236
rect 484032 7812 484084 7818
rect 484032 7754 484084 7760
rect 482284 3460 482336 3466
rect 482284 3402 482336 3408
rect 484044 480 484072 7754
rect 485228 3528 485280 3534
rect 485228 3470 485280 3476
rect 485240 480 485268 3470
rect 487632 480 487660 8230
rect 488828 480 488856 16546
rect 489012 3602 489040 499854
rect 489656 6322 489684 499854
rect 490300 233918 490328 499854
rect 491036 498166 491064 499854
rect 491588 499854 491662 499882
rect 492278 499882 492306 500140
rect 492922 499882 492950 500140
rect 493566 499882 493594 500140
rect 494210 499882 494238 500140
rect 494854 499882 494882 500140
rect 492278 499854 492352 499882
rect 491024 498160 491076 498166
rect 491024 498102 491076 498108
rect 490288 233912 490340 233918
rect 490288 233854 490340 233860
rect 489920 69080 489972 69086
rect 489920 69022 489972 69028
rect 489932 16574 489960 69022
rect 489932 16546 490696 16574
rect 489644 6316 489696 6322
rect 489644 6258 489696 6264
rect 489000 3596 489052 3602
rect 489000 3538 489052 3544
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 491588 6254 491616 499854
rect 492324 499574 492352 499854
rect 491956 499546 492352 499574
rect 491956 47598 491984 499546
rect 492324 499322 492352 499546
rect 492876 499854 492950 499882
rect 493520 499854 493594 499882
rect 494164 499854 494238 499882
rect 494808 499854 494882 499882
rect 495498 499882 495526 500140
rect 496142 499905 496170 500140
rect 496128 499896 496184 499905
rect 495498 499854 495572 499882
rect 492312 499316 492364 499322
rect 492312 499258 492364 499264
rect 492876 497554 492904 499854
rect 493520 497690 493548 499854
rect 493508 497684 493560 497690
rect 493508 497626 493560 497632
rect 492864 497548 492916 497554
rect 492864 497490 492916 497496
rect 493416 497480 493468 497486
rect 493416 497422 493468 497428
rect 493324 496868 493376 496874
rect 493324 496810 493376 496816
rect 491944 47592 491996 47598
rect 491944 47534 491996 47540
rect 493336 15910 493364 496810
rect 493428 26926 493456 497422
rect 494164 496874 494192 499854
rect 494808 497894 494836 499854
rect 494796 497888 494848 497894
rect 494796 497830 494848 497836
rect 494704 496936 494756 496942
rect 494704 496878 494756 496884
rect 494152 496868 494204 496874
rect 494152 496810 494204 496816
rect 493416 26920 493468 26926
rect 493416 26862 493468 26868
rect 493324 15904 493376 15910
rect 493324 15846 493376 15852
rect 494716 10334 494744 496878
rect 494808 14482 494836 497830
rect 495544 496194 495572 499854
rect 496786 499882 496814 500140
rect 497430 499882 497458 500140
rect 498074 499882 498102 500140
rect 498718 499882 498746 500140
rect 499362 499882 499390 500140
rect 500006 499882 500034 500140
rect 500650 499882 500678 500140
rect 501294 499882 501322 500140
rect 501938 499882 501966 500140
rect 502582 499882 502610 500140
rect 503226 499882 503254 500140
rect 503870 499882 503898 500140
rect 504514 499882 504542 500140
rect 505158 499882 505186 500140
rect 505802 499882 505830 500140
rect 506446 499882 506474 500140
rect 507090 499882 507118 500140
rect 507734 499882 507762 500140
rect 508378 499882 508406 500140
rect 509022 499882 509050 500140
rect 496128 499831 496184 499840
rect 496740 499854 496814 499882
rect 497384 499854 497458 499882
rect 498028 499854 498102 499882
rect 498672 499854 498746 499882
rect 499316 499854 499390 499882
rect 499960 499854 500034 499882
rect 500604 499854 500678 499882
rect 501248 499854 501322 499882
rect 501892 499854 501966 499882
rect 502536 499854 502610 499882
rect 503180 499854 503254 499882
rect 503824 499854 503898 499882
rect 504468 499854 504542 499882
rect 505112 499854 505186 499882
rect 505756 499854 505830 499882
rect 506400 499854 506474 499882
rect 507044 499854 507118 499882
rect 507688 499854 507762 499882
rect 508332 499854 508406 499882
rect 508976 499854 509050 499882
rect 509666 499882 509694 500140
rect 509666 499854 509740 499882
rect 496740 497962 496768 499854
rect 496728 497956 496780 497962
rect 496728 497898 496780 497904
rect 496176 497004 496228 497010
rect 496176 496946 496228 496952
rect 496084 496868 496136 496874
rect 496084 496810 496136 496816
rect 495532 496188 495584 496194
rect 495532 496130 495584 496136
rect 495438 39264 495494 39273
rect 495438 39199 495494 39208
rect 494796 14476 494848 14482
rect 494796 14418 494848 14424
rect 494704 10328 494756 10334
rect 494704 10270 494756 10276
rect 494704 9104 494756 9110
rect 494704 9046 494756 9052
rect 491576 6248 491628 6254
rect 491576 6190 491628 6196
rect 492310 4040 492366 4049
rect 492310 3975 492366 3984
rect 492324 480 492352 3975
rect 494716 480 494744 9046
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495452 354 495480 39199
rect 496096 19990 496124 496810
rect 496188 35290 496216 496946
rect 497384 482322 497412 499854
rect 498028 496942 498056 499854
rect 498016 496936 498068 496942
rect 498016 496878 498068 496884
rect 498672 496874 498700 499854
rect 499316 499390 499344 499854
rect 499304 499384 499356 499390
rect 499304 499326 499356 499332
rect 498660 496868 498712 496874
rect 498660 496810 498712 496816
rect 497372 482316 497424 482322
rect 497372 482258 497424 482264
rect 498200 352640 498252 352646
rect 498200 352582 498252 352588
rect 496176 35284 496228 35290
rect 496176 35226 496228 35232
rect 496084 19984 496136 19990
rect 496084 19926 496136 19932
rect 498212 3534 498240 352582
rect 498292 17332 498344 17338
rect 498292 17274 498344 17280
rect 498200 3528 498252 3534
rect 498200 3470 498252 3476
rect 498304 3346 498332 17274
rect 499960 6186 499988 499854
rect 500604 281518 500632 499854
rect 500592 281512 500644 281518
rect 500592 281454 500644 281460
rect 501248 33794 501276 499854
rect 501892 497010 501920 499854
rect 502536 498030 502564 499854
rect 503180 498098 503208 499854
rect 503168 498092 503220 498098
rect 503168 498034 503220 498040
rect 502524 498024 502576 498030
rect 502524 497966 502576 497972
rect 501880 497004 501932 497010
rect 501880 496946 501932 496952
rect 502340 496936 502392 496942
rect 502340 496878 502392 496884
rect 501236 33788 501288 33794
rect 501236 33730 501288 33736
rect 502352 16574 502380 496878
rect 503824 496874 503852 499854
rect 502984 496868 503036 496874
rect 502984 496810 503036 496816
rect 503812 496868 503864 496874
rect 503812 496810 503864 496816
rect 502996 29646 503024 496810
rect 502984 29640 503036 29646
rect 502984 29582 503036 29588
rect 504468 21486 504496 499854
rect 505112 106282 505140 499854
rect 505756 497622 505784 499854
rect 505744 497616 505796 497622
rect 505744 497558 505796 497564
rect 506400 480962 506428 499854
rect 507044 497486 507072 499854
rect 507032 497480 507084 497486
rect 507032 497422 507084 497428
rect 506388 480956 506440 480962
rect 506388 480898 506440 480904
rect 505100 106276 505152 106282
rect 505100 106218 505152 106224
rect 504456 21480 504508 21486
rect 504456 21422 504508 21428
rect 502352 16546 503024 16574
rect 499948 6180 500000 6186
rect 499948 6122 500000 6128
rect 499028 3528 499080 3534
rect 499028 3470 499080 3476
rect 498212 3318 498332 3346
rect 498212 480 498240 3318
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3470
rect 502996 480 503024 16546
rect 507688 4894 507716 499854
rect 508332 4962 508360 499854
rect 508504 498840 508556 498846
rect 508504 498782 508556 498788
rect 508320 4956 508372 4962
rect 508320 4898 508372 4904
rect 507676 4888 507728 4894
rect 507676 4830 507728 4836
rect 508516 3670 508544 498782
rect 508504 3664 508556 3670
rect 508504 3606 508556 3612
rect 508976 3194 509004 499854
rect 509712 496942 509740 499854
rect 509700 496936 509752 496942
rect 509700 496878 509752 496884
rect 509804 53106 509832 517919
rect 509896 224262 509924 522951
rect 510724 514321 510752 595410
rect 512092 569220 512144 569226
rect 512092 569162 512144 569168
rect 512000 555484 512052 555490
rect 512000 555426 512052 555432
rect 511170 529000 511226 529009
rect 511170 528935 511226 528944
rect 511078 526552 511134 526561
rect 511078 526487 511134 526496
rect 510986 520296 511042 520305
rect 510986 520231 511042 520240
rect 510802 519344 510858 519353
rect 510802 519279 510858 519288
rect 510710 514312 510766 514321
rect 510710 514247 510766 514256
rect 510816 514162 510844 519279
rect 511000 518894 511028 520231
rect 510632 514134 510844 514162
rect 510908 518866 511028 518894
rect 510066 513020 510122 513029
rect 510066 512955 510122 512964
rect 509974 511184 510030 511193
rect 509974 511119 510030 511128
rect 509884 224256 509936 224262
rect 509884 224198 509936 224204
rect 509792 53100 509844 53106
rect 509792 53042 509844 53048
rect 509988 8974 510016 511119
rect 510080 352646 510108 512955
rect 510434 510300 510490 510309
rect 510434 510235 510490 510244
rect 510250 505540 510306 505549
rect 510250 505475 510306 505484
rect 510264 497894 510292 505475
rect 510342 502140 510398 502149
rect 510342 502075 510398 502084
rect 510252 497888 510304 497894
rect 510252 497830 510304 497836
rect 510068 352640 510120 352646
rect 510068 352582 510120 352588
rect 510356 9042 510384 502075
rect 510448 493338 510476 510235
rect 510436 493332 510488 493338
rect 510436 493274 510488 493280
rect 510344 9036 510396 9042
rect 510344 8978 510396 8984
rect 509976 8968 510028 8974
rect 509976 8910 510028 8916
rect 510632 7614 510660 514134
rect 510908 514026 510936 518866
rect 510986 514448 511042 514457
rect 510986 514383 511042 514392
rect 510816 513998 510936 514026
rect 510710 507104 510766 507113
rect 510710 507039 510766 507048
rect 510724 500954 510752 507039
rect 510712 500948 510764 500954
rect 510712 500890 510764 500896
rect 510712 500812 510764 500818
rect 510712 500754 510764 500760
rect 510724 20670 510752 500754
rect 510816 220114 510844 513998
rect 511000 509234 511028 514383
rect 510908 509206 511028 509234
rect 510908 241466 510936 509206
rect 510986 505744 511042 505753
rect 510986 505679 511042 505688
rect 511000 500818 511028 505679
rect 510988 500812 511040 500818
rect 510988 500754 511040 500760
rect 510988 500676 511040 500682
rect 510988 500618 511040 500624
rect 511000 268394 511028 500618
rect 511092 349858 511120 526487
rect 511184 494834 511212 528935
rect 511262 507920 511318 507929
rect 511262 507855 511318 507864
rect 511276 500682 511304 507855
rect 511354 504384 511410 504393
rect 511354 504319 511410 504328
rect 511264 500676 511316 500682
rect 511264 500618 511316 500624
rect 511368 499322 511396 504319
rect 512012 503713 512040 555426
rect 511998 503704 512054 503713
rect 511998 503639 512054 503648
rect 511998 500984 512054 500993
rect 511998 500919 512054 500928
rect 511356 499316 511408 499322
rect 511356 499258 511408 499264
rect 512012 498846 512040 500919
rect 512104 500857 512132 569162
rect 512182 567896 512238 567905
rect 512182 567831 512238 567840
rect 512196 518265 512224 567831
rect 512276 558204 512328 558210
rect 512276 558146 512328 558152
rect 512288 526425 512316 558146
rect 513380 528896 513432 528902
rect 513380 528838 513432 528844
rect 513288 528624 513340 528630
rect 513286 528592 513288 528601
rect 513340 528592 513342 528601
rect 513286 528527 513342 528536
rect 512550 527232 512606 527241
rect 512550 527167 512606 527176
rect 512274 526416 512330 526425
rect 512274 526351 512330 526360
rect 512366 524512 512422 524521
rect 512366 524447 512422 524456
rect 512182 518256 512238 518265
rect 512182 518191 512238 518200
rect 512274 515672 512330 515681
rect 512274 515607 512330 515616
rect 512090 500848 512146 500857
rect 512090 500783 512146 500792
rect 512000 498840 512052 498846
rect 512000 498782 512052 498788
rect 511172 494828 511224 494834
rect 511172 494770 511224 494776
rect 511080 349852 511132 349858
rect 511080 349794 511132 349800
rect 510988 268388 511040 268394
rect 510988 268330 511040 268336
rect 510896 241460 510948 241466
rect 510896 241402 510948 241408
rect 510804 220108 510856 220114
rect 510804 220050 510856 220056
rect 512288 40730 512316 515607
rect 512380 225690 512408 524447
rect 512564 524362 512592 527167
rect 512642 524920 512698 524929
rect 512642 524855 512698 524864
rect 512656 524482 512684 524855
rect 512644 524476 512696 524482
rect 512644 524418 512696 524424
rect 512564 524334 512684 524362
rect 512550 523424 512606 523433
rect 512550 523359 512606 523368
rect 512458 522064 512514 522073
rect 512458 521999 512514 522008
rect 512472 281450 512500 521999
rect 512564 352578 512592 523359
rect 512656 493406 512684 524334
rect 512826 521792 512882 521801
rect 512826 521727 512882 521736
rect 512734 499896 512790 499905
rect 512734 499831 512790 499840
rect 512644 493400 512696 493406
rect 512644 493342 512696 493348
rect 512552 352572 512604 352578
rect 512552 352514 512604 352520
rect 512460 281444 512512 281450
rect 512460 281386 512512 281392
rect 512368 225684 512420 225690
rect 512368 225626 512420 225632
rect 512276 40724 512328 40730
rect 512276 40666 512328 40672
rect 510712 20664 510764 20670
rect 510712 20606 510764 20612
rect 510620 7608 510672 7614
rect 510620 7550 510672 7556
rect 512748 4826 512776 499831
rect 512840 7682 512868 521727
rect 512918 520704 512974 520713
rect 512918 520639 512974 520648
rect 512932 518894 512960 520639
rect 513286 519072 513342 519081
rect 513286 519007 513342 519016
rect 513300 518974 513328 519007
rect 513288 518968 513340 518974
rect 513288 518910 513340 518916
rect 512932 518866 513052 518894
rect 512918 506560 512974 506569
rect 512918 506495 512974 506504
rect 512932 494902 512960 506495
rect 512920 494896 512972 494902
rect 512920 494838 512972 494844
rect 513024 43450 513052 518866
rect 513194 516624 513250 516633
rect 513194 516559 513250 516568
rect 513208 516254 513236 516559
rect 513286 516352 513342 516361
rect 513286 516287 513342 516296
rect 513196 516248 513248 516254
rect 513196 516190 513248 516196
rect 513300 516186 513328 516287
rect 513288 516180 513340 516186
rect 513288 516122 513340 516128
rect 513196 516112 513248 516118
rect 513196 516054 513248 516060
rect 513208 515545 513236 516054
rect 513194 515536 513250 515545
rect 513194 515471 513250 515480
rect 513286 510776 513342 510785
rect 513286 510711 513342 510720
rect 513300 510678 513328 510711
rect 513288 510672 513340 510678
rect 513288 510614 513340 510620
rect 513286 509416 513342 509425
rect 513286 509351 513342 509360
rect 513300 509318 513328 509351
rect 513288 509312 513340 509318
rect 513288 509254 513340 509260
rect 513286 503976 513342 503985
rect 513286 503911 513342 503920
rect 513300 503742 513328 503911
rect 513288 503736 513340 503742
rect 513288 503678 513340 503684
rect 513286 502616 513342 502625
rect 513286 502551 513342 502560
rect 513300 502382 513328 502551
rect 513288 502376 513340 502382
rect 513288 502318 513340 502324
rect 513012 43444 513064 43450
rect 513012 43386 513064 43392
rect 512828 7676 512880 7682
rect 512828 7618 512880 7624
rect 512736 4820 512788 4826
rect 512736 4762 512788 4768
rect 510068 3460 510120 3466
rect 510068 3402 510120 3408
rect 506480 3188 506532 3194
rect 506480 3130 506532 3136
rect 508964 3188 509016 3194
rect 508964 3130 509016 3136
rect 506492 480 506520 3130
rect 510080 480 510108 3402
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 528838
rect 518164 528624 518216 528630
rect 518164 528566 518216 528572
rect 518176 431934 518204 528566
rect 520936 516118 520964 699654
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 525156 696992 525208 696998
rect 525156 696934 525208 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 521658 641744 521714 641753
rect 521658 641679 521714 641688
rect 521672 612377 521700 641679
rect 523684 641096 523736 641102
rect 523684 641038 523736 641044
rect 523696 632058 523724 641038
rect 523684 632052 523736 632058
rect 523684 631994 523736 632000
rect 521750 630728 521806 630737
rect 521750 630663 521806 630672
rect 521658 612368 521714 612377
rect 521658 612303 521714 612312
rect 520924 516112 520976 516118
rect 520924 516054 520976 516060
rect 521672 498166 521700 612303
rect 521764 598942 521792 630663
rect 521752 598936 521804 598942
rect 521752 598878 521804 598884
rect 525064 524476 525116 524482
rect 525064 524418 525116 524424
rect 522304 509312 522356 509318
rect 522304 509254 522356 509260
rect 521660 498160 521712 498166
rect 521660 498102 521712 498108
rect 518164 431928 518216 431934
rect 518164 431870 518216 431876
rect 516140 177404 516192 177410
rect 516140 177346 516192 177352
rect 516152 16574 516180 177346
rect 520280 177336 520332 177342
rect 520280 177278 520332 177284
rect 516152 16546 517192 16574
rect 517164 480 517192 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 177278
rect 522316 3534 522344 509254
rect 525076 3534 525104 524418
rect 525168 499458 525196 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 526444 643136 526496 643142
rect 526444 643078 526496 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 526456 533390 526484 643078
rect 530584 641028 530636 641034
rect 530584 640970 530636 640976
rect 526444 533384 526496 533390
rect 526444 533326 526496 533332
rect 527824 531616 527876 531622
rect 527824 531558 527876 531564
rect 526444 516248 526496 516254
rect 526444 516190 526496 516196
rect 525156 499452 525208 499458
rect 525156 499394 525208 499400
rect 526456 3602 526484 516190
rect 527836 16574 527864 531558
rect 530596 525774 530624 640970
rect 580172 632052 580224 632058
rect 580172 631994 580224 632000
rect 580184 630873 580212 631994
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 538864 616888 538916 616894
rect 538864 616830 538916 616836
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 538876 558278 538904 616830
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580262 578912 580318 578921
rect 580262 578847 580318 578856
rect 580172 578196 580224 578202
rect 580172 578138 580224 578144
rect 580184 577697 580212 578138
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 538864 558272 538916 558278
rect 538864 558214 538916 558220
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 549904 531752 549956 531758
rect 549904 531694 549956 531700
rect 534724 531548 534776 531554
rect 534724 531490 534776 531496
rect 530584 525768 530636 525774
rect 530584 525710 530636 525716
rect 531964 518968 532016 518974
rect 531964 518910 532016 518916
rect 530584 503736 530636 503742
rect 530584 503678 530636 503684
rect 527836 16546 527956 16574
rect 526444 3596 526496 3602
rect 526444 3538 526496 3544
rect 522304 3528 522356 3534
rect 522304 3470 522356 3476
rect 524236 3528 524288 3534
rect 524236 3470 524288 3476
rect 525064 3528 525116 3534
rect 525064 3470 525116 3476
rect 527824 3528 527876 3534
rect 527824 3470 527876 3476
rect 524248 480 524276 3470
rect 527836 480 527864 3470
rect 527928 3466 527956 16546
rect 530596 3670 530624 503678
rect 531976 3670 532004 518910
rect 530584 3664 530636 3670
rect 530584 3606 530636 3612
rect 531964 3664 532016 3670
rect 531964 3606 532016 3612
rect 531320 3596 531372 3602
rect 531320 3538 531372 3544
rect 527916 3460 527968 3466
rect 527916 3402 527968 3408
rect 531332 480 531360 3538
rect 534736 3534 534764 531490
rect 538864 531480 538916 531486
rect 538864 531422 538916 531428
rect 536104 516180 536156 516186
rect 536104 516122 536156 516128
rect 536116 153202 536144 516122
rect 536104 153196 536156 153202
rect 536104 153138 536156 153144
rect 538876 3738 538904 531422
rect 544384 510672 544436 510678
rect 544384 510614 544436 510620
rect 538864 3732 538916 3738
rect 538864 3674 538916 3680
rect 541992 3664 542044 3670
rect 541992 3606 542044 3612
rect 538404 3596 538456 3602
rect 538404 3538 538456 3544
rect 534724 3528 534776 3534
rect 534724 3470 534776 3476
rect 534908 3460 534960 3466
rect 534908 3402 534960 3408
rect 534920 480 534948 3402
rect 538416 480 538444 3538
rect 542004 480 542032 3606
rect 544396 3602 544424 510614
rect 545764 502376 545816 502382
rect 545764 502318 545816 502324
rect 544384 3596 544436 3602
rect 544384 3538 544436 3544
rect 545776 3466 545804 502318
rect 547880 496120 547932 496126
rect 547880 496062 547932 496068
rect 547892 16574 547920 496062
rect 547892 16546 548656 16574
rect 545488 3460 545540 3466
rect 545488 3402 545540 3408
rect 545764 3460 545816 3466
rect 545764 3402 545816 3408
rect 545500 480 545528 3402
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 549916 3534 549944 531694
rect 563060 530188 563112 530194
rect 563060 530130 563112 530136
rect 552664 496188 552716 496194
rect 552664 496130 552716 496136
rect 552020 354000 552072 354006
rect 552020 353942 552072 353948
rect 552032 16574 552060 353942
rect 552676 193186 552704 496130
rect 552664 193180 552716 193186
rect 552664 193122 552716 193128
rect 552032 16546 552704 16574
rect 549904 3528 549956 3534
rect 549904 3470 549956 3476
rect 552676 480 552704 16546
rect 559748 5024 559800 5030
rect 559748 4966 559800 4972
rect 556160 3732 556212 3738
rect 556160 3674 556212 3680
rect 556172 480 556200 3674
rect 559760 480 559788 4966
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563072 354 563100 530130
rect 565820 530052 565872 530058
rect 565820 529994 565872 530000
rect 565832 16574 565860 529994
rect 571984 529984 572036 529990
rect 571984 529926 572036 529932
rect 569960 527876 570012 527882
rect 569960 527818 570012 527824
rect 569972 16574 570000 527818
rect 571996 113150 572024 529926
rect 580172 525768 580224 525774
rect 580172 525710 580224 525716
rect 580184 524521 580212 525710
rect 580170 524512 580226 524521
rect 580170 524447 580226 524456
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580172 471980 580224 471986
rect 580172 471922 580224 471928
rect 580184 471481 580212 471922
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 579620 431928 579672 431934
rect 579620 431870 579672 431876
rect 579632 431633 579660 431870
rect 579618 431624 579674 431633
rect 579618 431559 579674 431568
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 578884 220856 578936 220862
rect 578884 220798 578936 220804
rect 571984 113144 572036 113150
rect 571984 113086 572036 113092
rect 565832 16546 566872 16574
rect 569972 16546 570368 16574
rect 566844 480 566872 16546
rect 570340 480 570368 16546
rect 573916 3596 573968 3602
rect 573916 3538 573968 3544
rect 573928 480 573956 3538
rect 578896 3534 578924 220798
rect 579896 219428 579948 219434
rect 579896 219370 579948 219376
rect 579908 219065 579936 219370
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579804 153196 579856 153202
rect 579804 153138 579856 153144
rect 579816 152697 579844 153138
rect 579802 152688 579858 152697
rect 579802 152623 579858 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580276 99521 580304 578847
rect 580354 564360 580410 564369
rect 580354 564295 580410 564304
rect 580368 554033 580396 564295
rect 580354 554024 580410 554033
rect 580354 553959 580410 553968
rect 582380 532024 582432 532030
rect 582380 531966 582432 531972
rect 580354 511320 580410 511329
rect 580354 511255 580410 511264
rect 580368 498710 580396 511255
rect 580356 498704 580408 498710
rect 580356 498646 580408 498652
rect 580448 489184 580500 489190
rect 580448 489126 580500 489132
rect 580356 486464 580408 486470
rect 580356 486406 580408 486412
rect 580368 378457 580396 486406
rect 580460 458153 580488 489126
rect 580446 458144 580502 458153
rect 580446 458079 580502 458088
rect 580354 378448 580410 378457
rect 580354 378383 580410 378392
rect 580356 341556 580408 341562
rect 580356 341498 580408 341504
rect 580368 325281 580396 341498
rect 580354 325272 580410 325281
rect 580354 325207 580410 325216
rect 580262 99512 580318 99521
rect 580262 99447 580318 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 582392 16574 582420 531966
rect 582392 16546 583432 16574
rect 581000 7744 581052 7750
rect 581000 7686 581052 7692
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 578884 3528 578936 3534
rect 578884 3470 578936 3476
rect 579804 3528 579856 3534
rect 579804 3470 579856 3476
rect 577412 3460 577464 3466
rect 577412 3402 577464 3408
rect 577424 480 577452 3402
rect 579816 480 579844 3470
rect 581012 480 581040 7686
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 583404 480 583432 16546
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3698 662632 3754 662688
rect 3514 662496 3570 662552
rect 3330 658144 3386 658200
rect 3790 553832 3846 553888
rect 3698 514800 3754 514856
rect 3606 501744 3662 501800
rect 3514 462576 3570 462632
rect 50986 663176 51042 663232
rect 46570 663040 46626 663096
rect 3422 449520 3478 449576
rect 46662 662904 46718 662960
rect 50066 661816 50122 661872
rect 49974 661680 50030 661736
rect 49330 661544 49386 661600
rect 48962 661408 49018 661464
rect 48870 661000 48926 661056
rect 48134 660592 48190 660648
rect 48042 660456 48098 660512
rect 47950 660320 48006 660376
rect 47950 421232 48006 421288
rect 48042 415384 48098 415440
rect 3146 410488 3202 410544
rect 48594 660184 48650 660240
rect 48134 409536 48190 409592
rect 48778 659912 48834 659968
rect 48594 584976 48650 585032
rect 48778 620064 48834 620120
rect 48686 579128 48742 579184
rect 48870 596672 48926 596728
rect 48962 590824 49018 590880
rect 49238 649304 49294 649360
rect 49146 631760 49202 631816
rect 49054 567432 49110 567488
rect 48778 555736 48834 555792
rect 49790 659640 49846 659696
rect 49606 655152 49662 655208
rect 50158 659776 50214 659832
rect 49606 643456 49662 643512
rect 50342 659640 50398 659696
rect 49422 637608 49478 637664
rect 49330 573280 49386 573336
rect 49238 561584 49294 561640
rect 49146 549888 49202 549944
rect 49422 544040 49478 544096
rect 49422 539552 49478 539608
rect 49422 538192 49478 538248
rect 49330 521600 49386 521656
rect 49330 520648 49386 520704
rect 49238 503104 49294 503160
rect 48870 496848 48926 496904
rect 48778 468016 48834 468072
rect 48318 444624 48374 444680
rect 48318 438812 48320 438832
rect 48320 438812 48372 438832
rect 48372 438812 48374 438832
rect 48318 438776 48374 438812
rect 48226 403688 48282 403744
rect 3422 397432 3478 397488
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 48318 392012 48374 392048
rect 48318 391992 48320 392012
rect 48320 391992 48372 392012
rect 48372 391992 48374 392012
rect 3514 306176 3570 306232
rect 3606 293120 3662 293176
rect 48318 386144 48374 386200
rect 48226 374448 48282 374504
rect 48134 368600 48190 368656
rect 48042 362752 48098 362808
rect 47950 351056 48006 351112
rect 47858 345208 47914 345264
rect 47950 281288 48006 281344
rect 47858 281152 47914 281208
rect 48134 280472 48190 280528
rect 48686 298424 48742 298480
rect 48778 292576 48834 292632
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 3146 136720 3202 136776
rect 3698 201864 3754 201920
rect 3606 188808 3662 188864
rect 3514 149776 3570 149832
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 19352 3478 19408
rect 4066 6432 4122 6488
rect 49606 497256 49662 497312
rect 49606 496848 49662 496904
rect 49514 491408 49570 491464
rect 48962 473864 49018 473920
rect 49146 432928 49202 432984
rect 49422 427080 49478 427136
rect 49422 380296 49478 380352
rect 49422 327664 49478 327720
rect 49330 321816 49386 321872
rect 49238 315968 49294 316024
rect 49146 304272 49202 304328
rect 49422 281016 49478 281072
rect 49330 280880 49386 280936
rect 49790 456356 49792 456376
rect 49792 456356 49844 456376
rect 49844 456356 49846 456376
rect 49790 456320 49846 456356
rect 50710 625912 50766 625968
rect 50986 532344 51042 532400
rect 50894 526496 50950 526552
rect 50802 508952 50858 509008
rect 50802 462168 50858 462224
rect 50710 456320 50766 456376
rect 51170 662768 51226 662824
rect 51262 659640 51318 659696
rect 51078 514800 51134 514856
rect 51262 485560 51318 485616
rect 51262 484336 51318 484392
rect 51262 450472 51318 450528
rect 52090 612720 52146 612776
rect 51998 607144 52054 607200
rect 51906 600752 51962 600808
rect 254582 658144 254638 658200
rect 254582 652296 254638 652352
rect 253938 646448 253994 646504
rect 254490 640600 254546 640656
rect 254398 634752 254454 634808
rect 254306 628904 254362 628960
rect 254030 623056 254086 623112
rect 254490 611380 254546 611416
rect 254490 611360 254492 611380
rect 254492 611360 254544 611380
rect 254544 611360 254546 611380
rect 254214 605512 254270 605568
rect 254122 599664 254178 599720
rect 254490 587988 254546 588024
rect 254490 587968 254492 587988
rect 254492 587968 254544 587988
rect 254544 587968 254546 587988
rect 253938 582120 253994 582176
rect 254490 576272 254546 576328
rect 253938 570424 253994 570480
rect 254674 617208 254730 617264
rect 254582 558728 254638 558784
rect 254398 552880 254454 552936
rect 254490 547032 254546 547088
rect 254766 593816 254822 593872
rect 254582 541204 254638 541240
rect 254582 541184 254584 541204
rect 254584 541184 254636 541204
rect 254636 541184 254638 541204
rect 254214 529488 254270 529544
rect 254030 523640 254086 523696
rect 254490 517792 254546 517848
rect 254398 511944 254454 512000
rect 254306 506096 254362 506152
rect 254214 500248 254270 500304
rect 254674 535336 254730 535392
rect 254582 494400 254638 494456
rect 51354 397840 51410 397896
rect 51354 356904 51410 356960
rect 51446 339360 51502 339416
rect 51354 281968 51410 282024
rect 51630 333512 51686 333568
rect 51538 310120 51594 310176
rect 51538 281832 51594 281888
rect 51446 280744 51502 280800
rect 51630 280608 51686 280664
rect 254398 482704 254454 482760
rect 254214 476856 254270 476912
rect 254490 471008 254546 471064
rect 254306 459312 254362 459368
rect 254398 441788 254454 441824
rect 254398 441768 254400 441788
rect 254400 441768 254452 441788
rect 254452 441768 254454 441788
rect 254214 430072 254270 430128
rect 254398 418376 254454 418432
rect 254306 406680 254362 406736
rect 254490 400832 254546 400888
rect 254490 395004 254546 395040
rect 254490 394984 254492 395004
rect 254492 394984 254544 395004
rect 254544 394984 254546 395004
rect 254490 389172 254492 389192
rect 254492 389172 254544 389192
rect 254544 389172 254546 389192
rect 254490 389136 254546 389172
rect 254214 383288 254270 383344
rect 254122 377440 254178 377496
rect 254398 371592 254454 371648
rect 254490 365764 254546 365800
rect 254490 365744 254492 365764
rect 254492 365744 254544 365764
rect 254544 365744 254546 365764
rect 253938 359896 253994 359952
rect 254490 354048 254546 354104
rect 253386 332016 253442 332072
rect 253202 331608 253258 331664
rect 52090 286456 52146 286512
rect 54574 278704 54630 278760
rect 59358 278024 59414 278080
rect 55862 223488 55918 223544
rect 57058 217368 57114 217424
rect 57150 209208 57206 209264
rect 57334 205128 57390 205184
rect 57334 201048 57390 201104
rect 57334 196968 57390 197024
rect 57242 192888 57298 192944
rect 57334 188808 57390 188864
rect 56690 184728 56746 184784
rect 56690 180648 56746 180704
rect 57334 176604 57336 176624
rect 57336 176604 57388 176624
rect 57388 176604 57390 176624
rect 57334 176568 57390 176604
rect 57242 172488 57298 172544
rect 57334 168408 57390 168464
rect 55862 164328 55918 164384
rect 57058 160248 57114 160304
rect 57058 156168 57114 156224
rect 57334 152088 57390 152144
rect 57334 148008 57390 148064
rect 57334 143928 57390 143984
rect 57426 139848 57482 139904
rect 57334 135768 57390 135824
rect 57518 123528 57574 123584
rect 57610 107208 57666 107264
rect 57702 103128 57758 103184
rect 57794 86808 57850 86864
rect 58898 127608 58954 127664
rect 58806 119448 58862 119504
rect 58990 111288 59046 111344
rect 59082 82728 59138 82784
rect 57886 78648 57942 78704
rect 59266 90888 59322 90944
rect 59450 276664 59506 276720
rect 59542 115368 59598 115424
rect 59450 94968 59506 95024
rect 59358 70488 59414 70544
rect 222842 215600 222898 215656
rect 60554 213832 60610 213888
rect 222290 212744 222346 212800
rect 223210 209888 223266 209944
rect 222934 207032 222990 207088
rect 222842 204176 222898 204232
rect 223026 201320 223082 201376
rect 222934 198464 222990 198520
rect 222842 189896 222898 189952
rect 222842 187040 222898 187096
rect 223486 195608 223542 195664
rect 223486 192752 223542 192808
rect 222290 184184 222346 184240
rect 223486 181328 223542 181384
rect 222658 178472 222714 178528
rect 222658 175616 222714 175672
rect 222382 172760 222438 172816
rect 222474 169904 222530 169960
rect 222934 167048 222990 167104
rect 223486 164192 223542 164248
rect 223026 161336 223082 161392
rect 222934 158480 222990 158536
rect 223486 155624 223542 155680
rect 222566 152768 222622 152824
rect 222474 144200 222530 144256
rect 223486 149912 223542 149968
rect 223486 147056 223542 147112
rect 223486 141344 223542 141400
rect 222934 138488 222990 138544
rect 222842 135632 222898 135688
rect 222474 132776 222530 132832
rect 223118 129920 223174 129976
rect 223486 127064 223542 127120
rect 222474 124208 222530 124264
rect 223210 121352 223266 121408
rect 223486 118496 223542 118552
rect 223486 115640 223542 115696
rect 222198 112784 222254 112840
rect 223486 109928 223542 109984
rect 222658 107072 222714 107128
rect 222842 104216 222898 104272
rect 223486 101360 223542 101416
rect 59818 99048 59874 99104
rect 223026 98504 223082 98560
rect 223118 95648 223174 95704
rect 223486 92792 223542 92848
rect 223486 89936 223542 89992
rect 223394 87080 223450 87136
rect 223486 84224 223542 84280
rect 223486 81388 223542 81424
rect 223486 81368 223488 81388
rect 223488 81368 223540 81388
rect 223540 81368 223542 81388
rect 222474 78548 222476 78568
rect 222476 78548 222528 78568
rect 222528 78548 222530 78568
rect 222474 78512 222530 78548
rect 222198 75692 222200 75712
rect 222200 75692 222252 75712
rect 222252 75692 222254 75712
rect 222198 75656 222254 75692
rect 59726 74568 59782 74624
rect 253570 331336 253626 331392
rect 254214 330656 254270 330712
rect 254490 324808 254546 324864
rect 254306 318960 254362 319016
rect 254214 307264 254270 307320
rect 254030 289720 254086 289776
rect 254306 283872 254362 283928
rect 254674 488572 254730 488608
rect 254674 488552 254676 488572
rect 254676 488552 254728 488572
rect 254728 488552 254730 488572
rect 254674 465160 254730 465216
rect 254674 453464 254730 453520
rect 254674 447616 254730 447672
rect 254674 435920 254730 435976
rect 254674 424224 254730 424280
rect 254674 412528 254730 412584
rect 254766 348200 254822 348256
rect 254674 342352 254730 342408
rect 254674 336504 254730 336560
rect 254674 313112 254730 313168
rect 254674 301416 254730 301472
rect 254674 295568 254730 295624
rect 222198 72800 222254 72856
rect 223486 69944 223542 70000
rect 223486 67088 223542 67144
rect 59634 66408 59690 66464
rect 257618 218592 257674 218648
rect 222842 64232 222898 64288
rect 59174 62328 59230 62384
rect 126978 61376 127034 61432
rect 74998 8880 75054 8936
rect 95790 10240 95846 10296
rect 136638 60016 136694 60072
rect 129738 59880 129794 59936
rect 147678 58520 147734 58576
rect 143538 10376 143594 10432
rect 165618 60152 165674 60208
rect 162490 3304 162546 3360
rect 187330 4800 187386 4856
rect 183742 3440 183798 3496
rect 278594 629992 278650 630048
rect 278686 610000 278742 610056
rect 296902 659776 296958 659832
rect 282734 641824 282790 641880
rect 304170 641688 304226 641744
rect 301962 640328 302018 640384
rect 306194 640464 306250 640520
rect 299110 639376 299166 639432
rect 282090 639240 282146 639296
rect 285402 639240 285458 639296
rect 288254 639240 288310 639296
rect 289634 639240 289690 639296
rect 298466 639240 298522 639296
rect 301962 600616 302018 600672
rect 280158 551248 280214 551304
rect 281630 573280 281686 573336
rect 287058 574640 287114 574696
rect 284298 571920 284354 571976
rect 282918 560904 282974 560960
rect 292670 574776 292726 574832
rect 294602 567976 294658 568032
rect 299478 582936 299534 582992
rect 299386 580216 299442 580272
rect 300674 598188 300730 598224
rect 300674 598168 300676 598188
rect 300676 598168 300728 598188
rect 300728 598168 300730 598188
rect 300674 581576 300730 581632
rect 302238 598848 302294 598904
rect 303434 600616 303490 600672
rect 306838 600616 306894 600672
rect 307574 600616 307630 600672
rect 302974 598848 303030 598904
rect 300950 592592 301006 592648
rect 296166 543360 296222 543416
rect 279790 542680 279846 542736
rect 292578 542680 292634 542736
rect 296166 542680 296222 542736
rect 297178 542408 297234 542464
rect 287886 539688 287942 539744
rect 298190 542816 298246 542872
rect 298926 542544 298982 542600
rect 299938 542408 299994 542464
rect 301870 543088 301926 543144
rect 283378 539552 283434 539608
rect 286138 539552 286194 539608
rect 287610 539552 287666 539608
rect 288622 539552 288678 539608
rect 289358 539552 289414 539608
rect 290554 539552 290610 539608
rect 290830 539552 290886 539608
rect 291566 539552 291622 539608
rect 293038 539552 293094 539608
rect 304078 542816 304134 542872
rect 304998 542680 305054 542736
rect 307022 543224 307078 543280
rect 306378 542408 306434 542464
rect 308494 542544 308550 542600
rect 308402 542408 308458 542464
rect 311898 568112 311954 568168
rect 309322 563760 309378 563816
rect 314658 558184 314714 558240
rect 312266 542816 312322 542872
rect 310702 542680 310758 542736
rect 309966 542544 310022 542600
rect 309414 542408 309470 542464
rect 311438 542408 311494 542464
rect 319626 598168 319682 598224
rect 319442 566344 319498 566400
rect 317510 543632 317566 543688
rect 320178 537308 320234 537364
rect 320362 512148 320418 512204
rect 320362 510824 320364 510844
rect 320364 510824 320416 510844
rect 320416 510824 320418 510844
rect 320362 510788 320418 510824
rect 320086 510108 320142 510164
rect 319350 509904 319406 509960
rect 320454 509496 320510 509552
rect 293222 332152 293278 332208
rect 293406 331472 293462 331528
rect 296074 498752 296130 498808
rect 295430 282104 295486 282160
rect 296534 331880 296590 331936
rect 296534 331744 296590 331800
rect 295982 204176 296038 204232
rect 297362 329704 297418 329760
rect 297270 324944 297326 325000
rect 297086 320184 297142 320240
rect 296994 301144 297050 301200
rect 296810 217640 296866 217696
rect 296810 202680 296866 202736
rect 296810 166776 296866 166832
rect 296810 157800 296866 157856
rect 296810 148824 296866 148880
rect 296810 135360 296866 135416
rect 296810 117408 296866 117464
rect 296994 102448 297050 102504
rect 297178 318824 297234 318880
rect 297454 328344 297510 328400
rect 297546 326304 297602 326360
rect 297730 323584 297786 323640
rect 297730 317464 297786 317520
rect 297730 316104 297786 316160
rect 297914 314744 297970 314800
rect 297914 312704 297970 312760
rect 298006 311344 298062 311400
rect 298006 306584 298062 306640
rect 298006 305224 298062 305280
rect 298650 308624 298706 308680
rect 298558 303864 298614 303920
rect 298006 302504 298062 302560
rect 297822 299104 297878 299160
rect 297730 296384 297786 296440
rect 297822 295024 297878 295080
rect 298006 291624 298062 291680
rect 297914 290264 297970 290320
rect 298006 288904 298062 288960
rect 298006 287544 298062 287600
rect 297638 284144 297694 284200
rect 297270 109928 297326 109984
rect 297454 218184 297510 218240
rect 297362 103944 297418 104000
rect 297546 192208 297602 192264
rect 297546 189216 297602 189272
rect 297546 142840 297602 142896
rect 297730 216144 297786 216200
rect 297730 214648 297786 214704
rect 297730 213152 297786 213208
rect 297730 211656 297786 211712
rect 297730 210160 297786 210216
rect 297730 208664 297786 208720
rect 297730 207168 297786 207224
rect 297730 205692 297786 205728
rect 297730 205672 297732 205692
rect 297732 205672 297784 205692
rect 297784 205672 297786 205692
rect 297730 201184 297786 201240
rect 297730 199688 297786 199744
rect 297730 198192 297786 198248
rect 297730 196696 297786 196752
rect 297730 195200 297786 195256
rect 297730 193704 297786 193760
rect 297730 190712 297786 190768
rect 297730 187720 297786 187776
rect 297730 186260 297732 186280
rect 297732 186260 297784 186280
rect 297784 186260 297786 186280
rect 297730 186224 297786 186260
rect 297730 184728 297786 184784
rect 297730 183232 297786 183288
rect 297730 181736 297786 181792
rect 297730 180240 297786 180296
rect 297730 178744 297786 178800
rect 297730 177248 297786 177304
rect 297730 175752 297786 175808
rect 297730 174256 297786 174312
rect 297730 172760 297786 172816
rect 297730 171264 297786 171320
rect 297730 169788 297786 169824
rect 297730 169768 297732 169788
rect 297732 169768 297784 169788
rect 297784 169768 297786 169788
rect 297730 168272 297786 168328
rect 297730 165280 297786 165336
rect 297730 163784 297786 163840
rect 297730 162288 297786 162344
rect 297730 160792 297786 160848
rect 297730 159296 297786 159352
rect 297730 156304 297786 156360
rect 297730 154808 297786 154864
rect 297730 153312 297786 153368
rect 297730 151836 297786 151872
rect 297730 151816 297732 151836
rect 297732 151816 297784 151836
rect 297784 151816 297786 151836
rect 297730 150320 297786 150376
rect 297730 147328 297786 147384
rect 297730 145832 297786 145888
rect 297730 144336 297786 144392
rect 297730 141344 297786 141400
rect 297730 139848 297786 139904
rect 297730 138352 297786 138408
rect 297730 136856 297786 136912
rect 297730 133864 297786 133920
rect 297730 132404 297732 132424
rect 297732 132404 297784 132424
rect 297784 132404 297786 132424
rect 297730 132368 297786 132404
rect 297730 130872 297786 130928
rect 297730 129376 297786 129432
rect 297730 127880 297786 127936
rect 297730 126384 297786 126440
rect 297730 124888 297786 124944
rect 297730 123392 297786 123448
rect 297730 121896 297786 121952
rect 297730 120400 297786 120456
rect 297730 118904 297786 118960
rect 297730 115912 297786 115968
rect 297730 114452 297732 114472
rect 297732 114452 297784 114472
rect 297784 114452 297786 114472
rect 297730 114416 297786 114452
rect 297730 112920 297786 112976
rect 297638 100952 297694 101008
rect 297454 99456 297510 99512
rect 297914 285504 297970 285560
rect 297914 106936 297970 106992
rect 297822 96464 297878 96520
rect 297086 91976 297142 92032
rect 299018 281288 299074 281344
rect 298834 97960 298890 98016
rect 298926 93472 298982 93528
rect 298006 90480 298062 90536
rect 299110 111424 299166 111480
rect 299202 108432 299258 108488
rect 299294 105440 299350 105496
rect 299662 322224 299718 322280
rect 299570 297744 299626 297800
rect 299570 282784 299626 282840
rect 299478 281424 299534 281480
rect 300674 331608 300730 331664
rect 305182 331200 305238 331256
rect 310334 332152 310390 332208
rect 319350 508292 319406 508328
rect 319350 508272 319352 508292
rect 319352 508272 319404 508292
rect 319404 508272 319406 508292
rect 320178 508068 320234 508124
rect 320086 506708 320142 506764
rect 319350 505572 319406 505608
rect 319350 505552 319352 505572
rect 319352 505552 319404 505572
rect 319404 505552 319406 505572
rect 320178 505348 320234 505404
rect 320086 504668 320142 504724
rect 319350 504192 319406 504248
rect 316130 331336 316186 331392
rect 320362 507388 320418 507444
rect 320546 508000 320602 508056
rect 320914 564984 320970 565040
rect 321006 555328 321062 555384
rect 322202 535336 322258 535392
rect 322202 532344 322258 532400
rect 321650 532208 321706 532264
rect 321558 527040 321614 527096
rect 322018 521872 322074 521928
rect 322018 520512 322074 520568
rect 321558 519308 321614 519344
rect 321558 519288 321560 519308
rect 321560 519288 321612 519308
rect 321612 519288 321614 519308
rect 321834 517792 321890 517848
rect 321558 517420 321560 517440
rect 321560 517420 321612 517440
rect 321612 517420 321614 517440
rect 321558 517384 321614 517420
rect 321834 515344 321890 515400
rect 321650 514120 321706 514176
rect 322110 514120 322166 514176
rect 320914 512080 320970 512136
rect 321558 511284 321614 511320
rect 321558 511264 321560 511284
rect 321560 511264 321612 511284
rect 321612 511264 321614 511284
rect 320914 340040 320970 340096
rect 321742 512624 321798 512680
rect 322110 512644 322166 512680
rect 322110 512624 322112 512644
rect 322112 512624 322164 512644
rect 322164 512624 322166 512644
rect 322478 536152 322534 536208
rect 322478 534384 322534 534440
rect 322386 533976 322442 534032
rect 322846 533296 322902 533352
rect 322478 531156 322480 531176
rect 322480 531156 322532 531176
rect 322532 531156 322534 531176
rect 322478 531120 322534 531156
rect 322386 530168 322442 530224
rect 322478 529760 322534 529816
rect 322754 528808 322810 528864
rect 322294 528400 322350 528456
rect 322478 528128 322534 528184
rect 322478 526768 322534 526824
rect 322478 525716 322480 525736
rect 322480 525716 322532 525736
rect 322532 525716 322534 525736
rect 322478 525680 322534 525716
rect 322570 524592 322626 524648
rect 322294 524456 322350 524512
rect 322478 523368 322534 523424
rect 322386 523096 322442 523152
rect 322478 522008 322534 522064
rect 322478 520648 322534 520704
rect 322478 517928 322534 517984
rect 322386 516332 322388 516352
rect 322388 516332 322440 516352
rect 322440 516332 322442 516352
rect 322386 516296 322442 516332
rect 322478 513440 322534 513496
rect 322846 519152 322902 519208
rect 322846 515480 322902 515536
rect 322386 504056 322442 504112
rect 322386 503376 322442 503432
rect 322386 502424 322442 502480
rect 321558 334600 321614 334656
rect 325698 518900 325754 518936
rect 325698 518880 325700 518900
rect 325700 518880 325752 518900
rect 325752 518880 325754 518900
rect 326986 518880 327042 518936
rect 327906 541048 327962 541104
rect 330482 530576 330538 530632
rect 332046 547032 332102 547088
rect 322938 331744 322994 331800
rect 350078 499296 350134 499352
rect 350078 498208 350134 498264
rect 349894 497528 349950 497584
rect 341890 332016 341946 332072
rect 348974 331472 349030 331528
rect 349986 326848 350042 326904
rect 350262 329024 350318 329080
rect 350170 327664 350226 327720
rect 350078 324944 350134 325000
rect 349802 315696 349858 315752
rect 349802 312160 349858 312216
rect 349986 305768 350042 305824
rect 349894 304408 349950 304464
rect 341062 147464 341118 147520
rect 340142 145288 340198 145344
rect 340050 138624 340106 138680
rect 299386 94968 299442 95024
rect 299018 88984 299074 89040
rect 296810 85992 296866 86048
rect 297178 77016 297234 77072
rect 296810 72528 296866 72584
rect 297178 68040 297234 68096
rect 298006 87488 298062 87544
rect 297546 84496 297602 84552
rect 297914 83000 297970 83056
rect 297914 81504 297970 81560
rect 298006 80028 298062 80064
rect 298006 80008 298008 80028
rect 298008 80008 298060 80028
rect 298060 80008 298062 80028
rect 297546 78512 297602 78568
rect 298006 75520 298062 75576
rect 298006 74024 298062 74080
rect 298006 69536 298062 69592
rect 297546 66544 297602 66600
rect 297362 65048 297418 65104
rect 297914 63552 297970 63608
rect 298006 62076 298062 62112
rect 298006 62056 298008 62076
rect 298008 62056 298060 62076
rect 298060 62056 298062 62076
rect 317418 60288 317474 60344
rect 297270 3576 297326 3632
rect 300766 3576 300822 3632
rect 340878 140936 340934 140992
rect 340234 119176 340290 119232
rect 340326 110472 340382 110528
rect 329194 3576 329250 3632
rect 340510 75656 340566 75712
rect 340970 114824 341026 114880
rect 342258 143112 342314 143168
rect 341246 132232 341302 132288
rect 341154 121352 341210 121408
rect 341338 112648 341394 112704
rect 341430 103944 341486 104000
rect 341522 101768 341578 101824
rect 341614 99592 341670 99648
rect 341706 97416 341762 97472
rect 342350 136584 342406 136640
rect 342442 134408 342498 134464
rect 342350 62600 342406 62656
rect 342534 130056 342590 130112
rect 342626 127880 342682 127936
rect 342534 80008 342590 80064
rect 342718 125704 342774 125760
rect 342810 123528 342866 123584
rect 342902 117000 342958 117056
rect 342902 108296 342958 108352
rect 342902 106120 342958 106176
rect 343086 93064 343142 93120
rect 342994 88712 343050 88768
rect 342902 86536 342958 86592
rect 343178 90888 343234 90944
rect 343086 79328 343142 79384
rect 343086 69128 343142 69184
rect 343178 66952 343234 67008
rect 343178 64776 343234 64832
rect 350722 301824 350778 301880
rect 350906 317464 350962 317520
rect 350906 307944 350962 308000
rect 350814 299104 350870 299160
rect 350722 291624 350778 291680
rect 350630 280744 350686 280800
rect 351090 288224 351146 288280
rect 350998 284144 351054 284200
rect 351458 497936 351514 497992
rect 351918 321544 351974 321600
rect 351458 314064 351514 314120
rect 351918 311344 351974 311400
rect 352010 306584 352066 306640
rect 351458 300464 351514 300520
rect 352102 297744 352158 297800
rect 351918 294344 351974 294400
rect 352102 292984 352158 293040
rect 351918 286864 351974 286920
rect 352378 318824 352434 318880
rect 352378 309984 352434 310040
rect 352286 290264 352342 290320
rect 352286 285504 352342 285560
rect 352470 296384 352526 296440
rect 353482 530576 353538 530632
rect 352746 323584 352802 323640
rect 352654 282784 352710 282840
rect 353482 291624 353538 291680
rect 355230 498888 355286 498944
rect 355506 497800 355562 497856
rect 355874 497392 355930 497448
rect 357162 550296 357218 550352
rect 357162 516160 357218 516216
rect 357162 499432 357218 499488
rect 357622 548528 357678 548584
rect 357438 547712 357494 547768
rect 357438 545944 357494 546000
rect 357438 544584 357494 544640
rect 357530 543496 357586 543552
rect 357438 539144 357494 539200
rect 357438 536732 357440 536752
rect 357440 536732 357492 536752
rect 357492 536732 357494 536752
rect 357438 536696 357494 536732
rect 357438 535372 357440 535392
rect 357440 535372 357492 535392
rect 357492 535372 357494 535392
rect 357438 535336 357494 535372
rect 357438 534928 357494 534984
rect 357530 534520 357586 534576
rect 357438 532344 357494 532400
rect 357530 531800 357586 531856
rect 357438 529488 357494 529544
rect 357438 526768 357494 526824
rect 357438 523640 357494 523696
rect 357714 533332 357716 533352
rect 357716 533332 357768 533352
rect 357768 533332 357770 533352
rect 357714 533296 357770 533332
rect 357438 519560 357494 519616
rect 357438 518744 357494 518800
rect 357530 517540 357586 517576
rect 357530 517520 357532 517540
rect 357532 517520 357584 517540
rect 357584 517520 357586 517540
rect 357438 517420 357440 517440
rect 357440 517420 357492 517440
rect 357492 517420 357494 517440
rect 357438 517384 357494 517420
rect 357438 514700 357440 514720
rect 357440 514700 357492 514720
rect 357492 514700 357494 514720
rect 357438 514664 357494 514700
rect 357438 512760 357494 512816
rect 357622 511536 357678 511592
rect 357438 511400 357494 511456
rect 357438 510312 357494 510368
rect 357438 508952 357494 509008
rect 357530 508680 357586 508736
rect 357438 507320 357494 507376
rect 357438 506232 357494 506288
rect 357530 505824 357586 505880
rect 357438 504600 357494 504656
rect 357438 503240 357494 503296
rect 357438 501880 357494 501936
rect 356886 497256 356942 497312
rect 357898 548392 357954 548448
rect 357990 543496 358046 543552
rect 357898 536560 357954 536616
rect 358450 540912 358506 540968
rect 358358 538056 358414 538112
rect 357898 526360 357954 526416
rect 358174 528536 358230 528592
rect 358082 525136 358138 525192
rect 357990 521872 358046 521928
rect 357806 510040 357862 510096
rect 357806 507728 357862 507784
rect 358266 519696 358322 519752
rect 358266 513168 358322 513224
rect 358542 527720 358598 527776
rect 358542 526904 358598 526960
rect 358450 522008 358506 522064
rect 358726 544992 358782 545048
rect 358818 543360 358874 543416
rect 358818 539280 358874 539336
rect 358634 525000 358690 525056
rect 358634 523776 358690 523832
rect 358542 516160 358598 516216
rect 358542 515072 358598 515128
rect 358726 503648 358782 503704
rect 358910 537784 358966 537840
rect 358910 532752 358966 532808
rect 359186 542272 359242 542328
rect 359094 521600 359150 521656
rect 401598 661272 401654 661328
rect 360934 641824 360990 641880
rect 365074 642232 365130 642288
rect 361946 639920 362002 639976
rect 365534 640056 365590 640112
rect 368938 641960 368994 642016
rect 369490 641688 369546 641744
rect 378046 640872 378102 640928
rect 390466 642096 390522 642152
rect 397090 641824 397146 641880
rect 398470 641688 398526 641744
rect 362590 639512 362646 639568
rect 362590 639376 362646 639432
rect 364062 639376 364118 639432
rect 381266 639512 381322 639568
rect 381358 639376 381414 639432
rect 381726 639396 381782 639432
rect 381726 639376 381728 639396
rect 381728 639376 381780 639396
rect 381780 639376 381782 639396
rect 385866 639396 385922 639432
rect 386142 639512 386198 639568
rect 385866 639376 385868 639396
rect 385868 639376 385920 639396
rect 385920 639376 385922 639396
rect 360934 551928 360990 551984
rect 361670 560224 361726 560280
rect 361762 558864 361818 558920
rect 361578 551792 361634 551848
rect 360842 550568 360898 550624
rect 363602 553424 363658 553480
rect 367282 598168 367338 598224
rect 368478 554240 368534 554296
rect 369030 552064 369086 552120
rect 370594 598304 370650 598360
rect 371146 598168 371202 598224
rect 369950 569200 370006 569256
rect 376114 597624 376170 597680
rect 376758 576816 376814 576872
rect 378322 583072 378378 583128
rect 378230 563896 378286 563952
rect 378874 598168 378930 598224
rect 379702 581848 379758 581904
rect 382462 581712 382518 581768
rect 382370 565120 382426 565176
rect 386602 580352 386658 580408
rect 388534 567976 388590 568032
rect 388442 560224 388498 560280
rect 389362 583752 389418 583808
rect 391202 596808 391258 596864
rect 392122 595448 392178 595504
rect 395526 586608 395582 586664
rect 396722 585656 396778 585712
rect 397458 550568 397514 550624
rect 398102 550568 398158 550624
rect 399574 559544 399630 559600
rect 359370 528264 359426 528320
rect 359278 520920 359334 520976
rect 359002 513304 359058 513360
rect 399942 546080 399998 546136
rect 400126 541524 400182 541580
rect 399850 536560 399906 536616
rect 399758 535608 399814 535664
rect 399758 533160 399814 533216
rect 399574 523640 399630 523696
rect 399482 507320 399538 507376
rect 400862 642232 400918 642288
rect 400494 561040 400550 561096
rect 400402 535404 400458 535460
rect 400310 525204 400366 525260
rect 400494 522960 400550 523016
rect 400770 538056 400826 538112
rect 400770 536288 400826 536344
rect 400678 527040 400734 527096
rect 400586 515480 400642 515536
rect 400218 504124 400274 504180
rect 399482 501608 399538 501664
rect 360658 499840 360714 499896
rect 360014 498072 360070 498128
rect 362590 499840 362646 499896
rect 361946 499160 362002 499216
rect 365166 499840 365222 499896
rect 365810 499432 365866 499488
rect 363878 497800 363934 497856
rect 364062 497800 364118 497856
rect 368386 499840 368442 499896
rect 367742 499432 367798 499488
rect 369674 499840 369730 499896
rect 370318 499840 370374 499896
rect 371606 498888 371662 498944
rect 369030 497936 369086 497992
rect 362958 497664 363014 497720
rect 364062 497392 364118 497448
rect 360842 497120 360898 497176
rect 374826 499840 374882 499896
rect 376114 499840 376170 499896
rect 376758 499840 376814 499896
rect 377402 499432 377458 499488
rect 376114 497392 376170 497448
rect 380622 499840 380678 499896
rect 381266 499840 381322 499896
rect 382554 499840 382610 499896
rect 382554 497528 382610 497584
rect 385130 499840 385186 499896
rect 385130 497800 385186 497856
rect 385774 497664 385830 497720
rect 387062 498072 387118 498128
rect 390282 499840 390338 499896
rect 387706 497936 387762 497992
rect 386418 497256 386474 497312
rect 391570 499704 391626 499760
rect 391570 497120 391626 497176
rect 392858 499840 392914 499896
rect 393502 499568 393558 499624
rect 395434 498072 395490 498128
rect 398654 499840 398710 499896
rect 400954 540640 401010 540696
rect 401690 551520 401746 551576
rect 401598 547440 401654 547496
rect 401690 544720 401746 544776
rect 401598 543088 401654 543144
rect 401598 541728 401654 541784
rect 401046 539280 401102 539336
rect 401598 536188 401600 536208
rect 401600 536188 401652 536208
rect 401652 536188 401654 536208
rect 401598 536152 401654 536188
rect 401966 540912 402022 540968
rect 401874 534656 401930 534712
rect 401874 533740 401876 533760
rect 401876 533740 401928 533760
rect 401928 533740 401930 533760
rect 401874 533704 401930 533740
rect 401782 533160 401838 533216
rect 401966 531800 402022 531856
rect 401966 530168 402022 530224
rect 401782 527040 401838 527096
rect 401598 520956 401600 520976
rect 401600 520956 401652 520976
rect 401652 520956 401654 520976
rect 401598 520920 401654 520956
rect 401598 520140 401600 520160
rect 401600 520140 401652 520160
rect 401652 520140 401654 520160
rect 401598 520104 401654 520140
rect 401598 516060 401600 516080
rect 401600 516060 401652 516080
rect 401652 516060 401654 516080
rect 401598 516024 401654 516060
rect 401598 513848 401654 513904
rect 401690 503240 401746 503296
rect 401966 527720 402022 527776
rect 402058 517384 402114 517440
rect 401966 515480 402022 515536
rect 401874 510448 401930 510504
rect 401874 508408 401930 508464
rect 401874 500248 401930 500304
rect 401782 499296 401838 499352
rect 402058 513440 402114 513496
rect 402242 526360 402298 526416
rect 402242 525000 402298 525056
rect 402426 532480 402482 532536
rect 403070 546352 403126 546408
rect 402886 530304 402942 530360
rect 402886 528944 402942 529000
rect 402886 528400 402942 528456
rect 403162 528808 403218 528864
rect 402886 524048 402942 524104
rect 402886 521736 402942 521792
rect 402518 518200 402574 518256
rect 402610 516180 402666 516216
rect 402610 516160 402612 516180
rect 402612 516160 402664 516180
rect 402664 516160 402666 516180
rect 402518 513204 402520 513224
rect 402520 513204 402572 513224
rect 402572 513204 402574 513224
rect 402518 513168 402574 513204
rect 402426 512760 402482 512816
rect 402334 511944 402390 512000
rect 402886 510720 402942 510776
rect 402886 509496 402942 509552
rect 402242 506404 402244 506424
rect 402244 506404 402296 506424
rect 402296 506404 402298 506424
rect 402242 506368 402298 506404
rect 402150 505960 402206 506016
rect 404910 509380 404966 509416
rect 404910 509360 404912 509380
rect 404912 509360 404964 509380
rect 404964 509360 404966 509380
rect 448610 177248 448666 177304
rect 474002 578992 474058 579048
rect 478694 636112 478750 636168
rect 478142 617752 478198 617808
rect 511998 661136 512054 661192
rect 484398 661000 484454 661056
rect 498198 661036 498200 661056
rect 498200 661036 498252 661056
rect 498252 661036 498254 661056
rect 498198 661000 498254 661036
rect 488538 660184 488594 660240
rect 500958 659776 501014 659832
rect 479706 596808 479762 596864
rect 477498 529624 477554 529680
rect 477498 528572 477500 528592
rect 477500 528572 477552 528592
rect 477552 528572 477554 528592
rect 477498 528536 477554 528572
rect 477498 527196 477554 527232
rect 477498 527176 477500 527196
rect 477500 527176 477552 527196
rect 477552 527176 477554 527196
rect 481822 532616 481878 532672
rect 482926 529896 482982 529952
rect 484674 532616 484730 532672
rect 488998 532616 489054 532672
rect 501878 532616 501934 532672
rect 500958 532480 501014 532536
rect 489550 529488 489606 529544
rect 502430 529488 502486 529544
rect 504178 529488 504234 529544
rect 479154 527448 479210 527504
rect 479062 526088 479118 526144
rect 477498 525836 477554 525872
rect 477498 525816 477500 525836
rect 477500 525816 477552 525836
rect 477552 525816 477554 525836
rect 477958 525580 477960 525600
rect 477960 525580 478012 525600
rect 478012 525580 478014 525600
rect 477958 525544 478014 525580
rect 478694 525000 478750 525056
rect 477498 523368 477554 523424
rect 477498 523096 477554 523152
rect 478418 522008 478474 522064
rect 477958 521736 478014 521792
rect 477498 520648 477554 520704
rect 477590 517928 477646 517984
rect 477498 517656 477554 517712
rect 477590 513848 477646 513904
rect 477498 513440 477554 513496
rect 477590 512760 477646 512816
rect 477590 511128 477646 511184
rect 477866 510584 477922 510640
rect 477498 510448 477554 510504
rect 477498 509360 477554 509416
rect 477498 505688 477554 505744
rect 477498 505280 477554 505336
rect 477590 504328 477646 504384
rect 477498 503920 477554 503976
rect 477498 502560 477554 502616
rect 477498 501608 477554 501664
rect 477498 500112 477554 500168
rect 478234 516976 478290 517032
rect 478142 507048 478198 507104
rect 478602 520240 478658 520296
rect 478510 519288 478566 519344
rect 478510 516840 478566 516896
rect 478510 507864 478566 507920
rect 478694 519016 478750 519072
rect 478970 515208 479026 515264
rect 478786 512896 478842 512952
rect 478786 508272 478842 508328
rect 478786 500928 478842 500984
rect 510618 526496 510674 526552
rect 509882 522960 509938 523016
rect 509790 517928 509846 517984
rect 479246 514800 479302 514856
rect 479430 506504 479486 506560
rect 479338 502968 479394 503024
rect 496128 499840 496184 499896
rect 495438 39208 495494 39264
rect 492310 3984 492366 4040
rect 511170 528944 511226 529000
rect 511078 526496 511134 526552
rect 510986 520240 511042 520296
rect 510802 519288 510858 519344
rect 510710 514256 510766 514312
rect 510066 512964 510122 513020
rect 509974 511128 510030 511184
rect 510434 510244 510490 510300
rect 510250 505484 510306 505540
rect 510342 502084 510398 502140
rect 510986 514392 511042 514448
rect 510710 507048 510766 507104
rect 510986 505688 511042 505744
rect 511262 507864 511318 507920
rect 511354 504328 511410 504384
rect 511998 503648 512054 503704
rect 511998 500928 512054 500984
rect 512182 567840 512238 567896
rect 513286 528572 513288 528592
rect 513288 528572 513340 528592
rect 513340 528572 513342 528592
rect 513286 528536 513342 528572
rect 512550 527176 512606 527232
rect 512274 526360 512330 526416
rect 512366 524456 512422 524512
rect 512182 518200 512238 518256
rect 512274 515616 512330 515672
rect 512090 500792 512146 500848
rect 512642 524864 512698 524920
rect 512550 523368 512606 523424
rect 512458 522008 512514 522064
rect 512826 521736 512882 521792
rect 512734 499840 512790 499896
rect 512918 520648 512974 520704
rect 513286 519016 513342 519072
rect 512918 506504 512974 506560
rect 513194 516568 513250 516624
rect 513286 516296 513342 516352
rect 513194 515480 513250 515536
rect 513286 510720 513342 510776
rect 513286 509360 513342 509416
rect 513286 503920 513342 503976
rect 513286 502560 513342 502616
rect 580170 697176 580226 697232
rect 521658 641688 521714 641744
rect 521750 630672 521806 630728
rect 521658 612312 521714 612368
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580262 578856 580318 578912
rect 580170 577632 580226 577688
rect 579894 537784 579950 537840
rect 580170 524456 580226 524512
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 579618 431568 579674 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 580170 312024 580226 312080
rect 579618 298696 579674 298752
rect 579894 272176 579950 272232
rect 579802 258848 579858 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 579894 219000 579950 219056
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 580170 165824 580226 165880
rect 579802 152632 579858 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 580170 112784 580226 112840
rect 580354 564304 580410 564360
rect 580354 553968 580410 554024
rect 580354 511264 580410 511320
rect 580446 458088 580502 458144
rect 580354 378392 580410 378448
rect 580354 325216 580410 325272
rect 580262 99456 580318 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684164 480 684404
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect -960 671198 674 671258
rect -960 671122 480 671198
rect 614 671122 674 671198
rect -960 671108 674 671122
rect 246 671062 674 671108
rect 246 670714 306 671062
rect 279366 670714 279372 670716
rect 246 670654 279372 670714
rect 279366 670652 279372 670654
rect 279436 670652 279442 670716
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect 50981 663234 51047 663237
rect 283414 663234 283420 663236
rect 50981 663232 283420 663234
rect 50981 663176 50986 663232
rect 51042 663176 283420 663232
rect 50981 663174 283420 663176
rect 50981 663171 51047 663174
rect 283414 663172 283420 663174
rect 283484 663172 283490 663236
rect 46565 663098 46631 663101
rect 286174 663098 286180 663100
rect 46565 663096 286180 663098
rect 46565 663040 46570 663096
rect 46626 663040 286180 663096
rect 46565 663038 286180 663040
rect 46565 663035 46631 663038
rect 286174 663036 286180 663038
rect 286244 663036 286250 663100
rect 46657 662962 46723 662965
rect 317638 662962 317644 662964
rect 46657 662960 317644 662962
rect 46657 662904 46662 662960
rect 46718 662904 317644 662960
rect 46657 662902 317644 662904
rect 46657 662899 46723 662902
rect 317638 662900 317644 662902
rect 317708 662900 317714 662964
rect 51165 662826 51231 662829
rect 403014 662826 403020 662828
rect 51165 662824 403020 662826
rect 51165 662768 51170 662824
rect 51226 662768 403020 662824
rect 51165 662766 403020 662768
rect 51165 662763 51231 662766
rect 403014 662764 403020 662766
rect 403084 662764 403090 662828
rect 3693 662690 3759 662693
rect 481582 662690 481588 662692
rect 3693 662688 481588 662690
rect 3693 662632 3698 662688
rect 3754 662632 481588 662688
rect 3693 662630 481588 662632
rect 3693 662627 3759 662630
rect 481582 662628 481588 662630
rect 481652 662628 481658 662692
rect 3509 662554 3575 662557
rect 495382 662554 495388 662556
rect 3509 662552 495388 662554
rect 3509 662496 3514 662552
rect 3570 662496 495388 662552
rect 3509 662494 495388 662496
rect 3509 662491 3575 662494
rect 495382 662492 495388 662494
rect 495452 662492 495458 662556
rect 50061 661874 50127 661877
rect 290958 661874 290964 661876
rect 50061 661872 290964 661874
rect 50061 661816 50066 661872
rect 50122 661816 290964 661872
rect 50061 661814 290964 661816
rect 50061 661811 50127 661814
rect 290958 661812 290964 661814
rect 291028 661812 291034 661876
rect 49969 661738 50035 661741
rect 295926 661738 295932 661740
rect 49969 661736 295932 661738
rect 49969 661680 49974 661736
rect 50030 661680 295932 661736
rect 49969 661678 295932 661680
rect 49969 661675 50035 661678
rect 295926 661676 295932 661678
rect 295996 661676 296002 661740
rect 49325 661602 49391 661605
rect 304206 661602 304212 661604
rect 49325 661600 304212 661602
rect 49325 661544 49330 661600
rect 49386 661544 304212 661600
rect 49325 661542 304212 661544
rect 49325 661539 49391 661542
rect 304206 661540 304212 661542
rect 304276 661540 304282 661604
rect 48957 661466 49023 661469
rect 305494 661466 305500 661468
rect 48957 661464 305500 661466
rect 48957 661408 48962 661464
rect 49018 661408 305500 661464
rect 48957 661406 305500 661408
rect 48957 661403 49023 661406
rect 305494 661404 305500 661406
rect 305564 661404 305570 661468
rect 401593 661332 401659 661333
rect 49366 661268 49372 661332
rect 49436 661330 49442 661332
rect 308622 661330 308628 661332
rect 49436 661270 308628 661330
rect 49436 661268 49442 661270
rect 308622 661268 308628 661270
rect 308692 661268 308698 661332
rect 401542 661268 401548 661332
rect 401612 661330 401659 661332
rect 401612 661328 401704 661330
rect 401654 661272 401704 661328
rect 401612 661270 401704 661272
rect 401612 661268 401659 661270
rect 401593 661267 401659 661268
rect 49550 661132 49556 661196
rect 49620 661194 49626 661196
rect 309358 661194 309364 661196
rect 49620 661134 309364 661194
rect 49620 661132 49626 661134
rect 309358 661132 309364 661134
rect 309428 661132 309434 661196
rect 511993 661194 512059 661197
rect 512126 661194 512132 661196
rect 511993 661192 512132 661194
rect 511993 661136 511998 661192
rect 512054 661136 512132 661192
rect 511993 661134 512132 661136
rect 511993 661131 512059 661134
rect 512126 661132 512132 661134
rect 512196 661132 512202 661196
rect 48865 661058 48931 661061
rect 309174 661058 309180 661060
rect 48865 661056 309180 661058
rect 48865 661000 48870 661056
rect 48926 661000 309180 661056
rect 48865 660998 309180 661000
rect 48865 660995 48931 660998
rect 309174 660996 309180 660998
rect 309244 660996 309250 661060
rect 484393 661058 484459 661061
rect 484894 661058 484900 661060
rect 484393 661056 484900 661058
rect 484393 661000 484398 661056
rect 484454 661000 484900 661056
rect 484393 660998 484900 661000
rect 484393 660995 484459 660998
rect 484894 660996 484900 660998
rect 484964 660996 484970 661060
rect 498193 661058 498259 661061
rect 499430 661058 499436 661060
rect 498193 661056 499436 661058
rect 498193 661000 498198 661056
rect 498254 661000 499436 661056
rect 498193 660998 499436 661000
rect 498193 660995 498259 660998
rect 499430 660996 499436 660998
rect 499500 660996 499506 661060
rect 48129 660650 48195 660653
rect 291694 660650 291700 660652
rect 48129 660648 291700 660650
rect 48129 660592 48134 660648
rect 48190 660592 291700 660648
rect 48129 660590 291700 660592
rect 48129 660587 48195 660590
rect 291694 660588 291700 660590
rect 291764 660588 291770 660652
rect 48037 660514 48103 660517
rect 295006 660514 295012 660516
rect 48037 660512 295012 660514
rect 48037 660456 48042 660512
rect 48098 660456 295012 660512
rect 48037 660454 295012 660456
rect 48037 660451 48103 660454
rect 295006 660452 295012 660454
rect 295076 660452 295082 660516
rect 47945 660378 48011 660381
rect 299974 660378 299980 660380
rect 47945 660376 299980 660378
rect 47945 660320 47950 660376
rect 48006 660320 299980 660376
rect 47945 660318 299980 660320
rect 47945 660315 48011 660318
rect 299974 660316 299980 660318
rect 300044 660316 300050 660380
rect 48589 660242 48655 660245
rect 308806 660242 308812 660244
rect 48589 660240 308812 660242
rect 48589 660184 48594 660240
rect 48650 660184 308812 660240
rect 48589 660182 308812 660184
rect 48589 660179 48655 660182
rect 308806 660180 308812 660182
rect 308876 660180 308882 660244
rect 488533 660242 488599 660245
rect 489126 660242 489132 660244
rect 488533 660240 489132 660242
rect 488533 660184 488538 660240
rect 488594 660184 489132 660240
rect 488533 660182 489132 660184
rect 488533 660179 488599 660182
rect 489126 660180 489132 660182
rect 489196 660180 489202 660244
rect 49182 660044 49188 660108
rect 49252 660106 49258 660108
rect 310462 660106 310468 660108
rect 49252 660046 310468 660106
rect 49252 660044 49258 660046
rect 310462 660044 310468 660046
rect 310532 660044 310538 660108
rect 48773 659970 48839 659973
rect 311934 659970 311940 659972
rect 48773 659968 311940 659970
rect 48773 659912 48778 659968
rect 48834 659912 311940 659968
rect 48773 659910 311940 659912
rect 48773 659907 48839 659910
rect 311934 659908 311940 659910
rect 312004 659908 312010 659972
rect 50153 659836 50219 659837
rect 50102 659834 50108 659836
rect 50062 659774 50108 659834
rect 50172 659832 50219 659836
rect 50214 659776 50219 659832
rect 50102 659772 50108 659774
rect 50172 659772 50219 659776
rect 50153 659771 50219 659772
rect 296897 659834 296963 659837
rect 297214 659834 297220 659836
rect 296897 659832 297220 659834
rect 296897 659776 296902 659832
rect 296958 659776 297220 659832
rect 296897 659774 297220 659776
rect 296897 659771 296963 659774
rect 297214 659772 297220 659774
rect 297284 659772 297290 659836
rect 500953 659834 501019 659837
rect 502006 659834 502012 659836
rect 500953 659832 502012 659834
rect 500953 659776 500958 659832
rect 501014 659776 502012 659832
rect 500953 659774 502012 659776
rect 500953 659771 501019 659774
rect 502006 659772 502012 659774
rect 502076 659772 502082 659836
rect 49785 659700 49851 659701
rect 49734 659698 49740 659700
rect 49694 659638 49740 659698
rect 49804 659696 49851 659700
rect 49846 659640 49851 659696
rect 49734 659636 49740 659638
rect 49804 659636 49851 659640
rect 49918 659636 49924 659700
rect 49988 659698 49994 659700
rect 50337 659698 50403 659701
rect 51257 659700 51323 659701
rect 51206 659698 51212 659700
rect 49988 659696 50403 659698
rect 49988 659640 50342 659696
rect 50398 659640 50403 659696
rect 49988 659638 50403 659640
rect 51166 659638 51212 659698
rect 51276 659696 51323 659700
rect 51318 659640 51323 659696
rect 49988 659636 49994 659638
rect 49785 659635 49851 659636
rect 50337 659635 50403 659638
rect 51206 659636 51212 659638
rect 51276 659636 51323 659640
rect 51257 659635 51323 659636
rect -960 658202 480 658292
rect 3325 658202 3391 658205
rect 254577 658202 254643 658205
rect -960 658200 3391 658202
rect -960 658144 3330 658200
rect 3386 658144 3391 658200
rect -960 658142 3391 658144
rect 251804 658200 254643 658202
rect 251804 658144 254582 658200
rect 254638 658144 254643 658200
rect 251804 658142 254643 658144
rect -960 658052 480 658142
rect 3325 658139 3391 658142
rect 254577 658139 254643 658142
rect 583520 657236 584960 657476
rect 49601 655210 49667 655213
rect 49601 655208 52164 655210
rect 49601 655152 49606 655208
rect 49662 655152 52164 655208
rect 49601 655150 52164 655152
rect 49601 655147 49667 655150
rect 254577 652354 254643 652357
rect 251804 652352 254643 652354
rect 251804 652296 254582 652352
rect 254638 652296 254643 652352
rect 251804 652294 254643 652296
rect 254577 652291 254643 652294
rect 49233 649362 49299 649365
rect 49233 649360 52164 649362
rect 49233 649304 49238 649360
rect 49294 649304 52164 649360
rect 49233 649302 52164 649304
rect 49233 649299 49299 649302
rect 253933 646506 253999 646509
rect 251804 646504 253999 646506
rect 251804 646448 253938 646504
rect 253994 646448 253999 646504
rect 251804 646446 253999 646448
rect 253933 646443 253999 646446
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 49601 643514 49667 643517
rect 49601 643512 52164 643514
rect 49601 643456 49606 643512
rect 49662 643456 52164 643512
rect 49601 643454 52164 643456
rect 49601 643451 49667 643454
rect 365069 642290 365135 642293
rect 400857 642290 400923 642293
rect 365069 642288 400923 642290
rect 365069 642232 365074 642288
rect 365130 642232 400862 642288
rect 400918 642232 400923 642288
rect 365069 642230 400923 642232
rect 365069 642227 365135 642230
rect 400857 642227 400923 642230
rect 359406 642092 359412 642156
rect 359476 642154 359482 642156
rect 390461 642154 390527 642157
rect 359476 642152 390527 642154
rect 359476 642096 390466 642152
rect 390522 642096 390527 642152
rect 359476 642094 390527 642096
rect 359476 642092 359482 642094
rect 390461 642091 390527 642094
rect 368933 642018 368999 642021
rect 398598 642018 398604 642020
rect 368933 642016 398604 642018
rect 368933 641960 368938 642016
rect 368994 641960 398604 642016
rect 368933 641958 398604 641960
rect 368933 641955 368999 641958
rect 398598 641956 398604 641958
rect 398668 641956 398674 642020
rect 282729 641882 282795 641885
rect 293166 641882 293172 641884
rect 282729 641880 293172 641882
rect 282729 641824 282734 641880
rect 282790 641824 293172 641880
rect 282729 641822 293172 641824
rect 282729 641819 282795 641822
rect 293166 641820 293172 641822
rect 293236 641820 293242 641884
rect 360929 641882 360995 641885
rect 397085 641882 397151 641885
rect 360929 641880 397151 641882
rect 360929 641824 360934 641880
rect 360990 641824 397090 641880
rect 397146 641824 397151 641880
rect 360929 641822 397151 641824
rect 360929 641819 360995 641822
rect 397085 641819 397151 641822
rect 304165 641746 304231 641749
rect 311014 641746 311020 641748
rect 304165 641744 311020 641746
rect 304165 641688 304170 641744
rect 304226 641688 311020 641744
rect 304165 641686 311020 641688
rect 304165 641683 304231 641686
rect 311014 641684 311020 641686
rect 311084 641684 311090 641748
rect 363454 641684 363460 641748
rect 363524 641746 363530 641748
rect 369485 641746 369551 641749
rect 363524 641744 369551 641746
rect 363524 641688 369490 641744
rect 369546 641688 369551 641744
rect 363524 641686 369551 641688
rect 363524 641684 363530 641686
rect 369485 641683 369551 641686
rect 398465 641746 398531 641749
rect 521653 641746 521719 641749
rect 398465 641744 521719 641746
rect 398465 641688 398470 641744
rect 398526 641688 521658 641744
rect 521714 641688 521719 641744
rect 398465 641686 521719 641688
rect 398465 641683 398531 641686
rect 521653 641683 521719 641686
rect 307518 640868 307524 640932
rect 307588 640930 307594 640932
rect 378041 640930 378107 640933
rect 307588 640928 378107 640930
rect 307588 640872 378046 640928
rect 378102 640872 378107 640928
rect 307588 640870 378107 640872
rect 307588 640868 307594 640870
rect 378041 640867 378107 640870
rect 254485 640658 254551 640661
rect 251804 640656 254551 640658
rect 251804 640600 254490 640656
rect 254546 640600 254551 640656
rect 251804 640598 254551 640600
rect 254485 640595 254551 640598
rect 306189 640522 306255 640525
rect 355358 640522 355364 640524
rect 306189 640520 355364 640522
rect 306189 640464 306194 640520
rect 306250 640464 355364 640520
rect 306189 640462 355364 640464
rect 306189 640459 306255 640462
rect 355358 640460 355364 640462
rect 355428 640460 355434 640524
rect 301957 640386 302023 640389
rect 355174 640386 355180 640388
rect 301957 640384 355180 640386
rect 301957 640328 301962 640384
rect 302018 640328 355180 640384
rect 301957 640326 355180 640328
rect 301957 640323 302023 640326
rect 355174 640324 355180 640326
rect 355244 640324 355250 640388
rect 365529 640114 365595 640117
rect 354630 640112 365595 640114
rect 354630 640056 365534 640112
rect 365590 640056 365595 640112
rect 354630 640054 365595 640056
rect 303470 639508 303476 639572
rect 303540 639570 303546 639572
rect 354630 639570 354690 640054
rect 365529 640051 365595 640054
rect 361941 639978 362007 639981
rect 362534 639978 362540 639980
rect 361941 639976 362540 639978
rect 361941 639920 361946 639976
rect 362002 639920 362540 639976
rect 361941 639918 362540 639920
rect 361941 639915 362007 639918
rect 362534 639916 362540 639918
rect 362604 639916 362610 639980
rect 303540 639510 354690 639570
rect 303540 639508 303546 639510
rect 362350 639508 362356 639572
rect 362420 639570 362426 639572
rect 362585 639570 362651 639573
rect 362420 639568 362651 639570
rect 362420 639512 362590 639568
rect 362646 639512 362651 639568
rect 362420 639510 362651 639512
rect 362420 639508 362426 639510
rect 362585 639507 362651 639510
rect 381261 639570 381327 639573
rect 386137 639570 386203 639573
rect 381261 639568 386203 639570
rect 381261 639512 381266 639568
rect 381322 639512 386142 639568
rect 386198 639512 386203 639568
rect 381261 639510 386203 639512
rect 381261 639507 381327 639510
rect 386137 639507 386203 639510
rect 298318 639372 298324 639436
rect 298388 639434 298394 639436
rect 299105 639434 299171 639437
rect 298388 639432 299171 639434
rect 298388 639376 299110 639432
rect 299166 639376 299171 639432
rect 298388 639374 299171 639376
rect 298388 639372 298394 639374
rect 299105 639371 299171 639374
rect 362585 639434 362651 639437
rect 364057 639436 364123 639437
rect 362718 639434 362724 639436
rect 362585 639432 362724 639434
rect 362585 639376 362590 639432
rect 362646 639376 362724 639432
rect 362585 639374 362724 639376
rect 362585 639371 362651 639374
rect 362718 639372 362724 639374
rect 362788 639372 362794 639436
rect 364006 639434 364012 639436
rect 363966 639374 364012 639434
rect 364076 639432 364123 639436
rect 381353 639434 381419 639437
rect 364118 639376 364123 639432
rect 364006 639372 364012 639374
rect 364076 639372 364123 639376
rect 364057 639371 364123 639372
rect 373950 639432 381419 639434
rect 373950 639376 381358 639432
rect 381414 639376 381419 639432
rect 373950 639374 381419 639376
rect 282085 639298 282151 639301
rect 285397 639300 285463 639301
rect 288249 639300 288315 639301
rect 282678 639298 282684 639300
rect 282085 639296 282684 639298
rect 282085 639240 282090 639296
rect 282146 639240 282684 639296
rect 282085 639238 282684 639240
rect 282085 639235 282151 639238
rect 282678 639236 282684 639238
rect 282748 639236 282754 639300
rect 285397 639296 285444 639300
rect 285508 639298 285514 639300
rect 288198 639298 288204 639300
rect 285397 639240 285402 639296
rect 285397 639236 285444 639240
rect 285508 639238 285554 639298
rect 288158 639238 288204 639298
rect 288268 639296 288315 639300
rect 288310 639240 288315 639296
rect 285508 639236 285514 639238
rect 288198 639236 288204 639238
rect 288268 639236 288315 639240
rect 289486 639236 289492 639300
rect 289556 639298 289562 639300
rect 289629 639298 289695 639301
rect 289556 639296 289695 639298
rect 289556 639240 289634 639296
rect 289690 639240 289695 639296
rect 289556 639238 289695 639240
rect 289556 639236 289562 639238
rect 285397 639235 285463 639236
rect 288249 639235 288315 639236
rect 289629 639235 289695 639238
rect 298461 639300 298527 639301
rect 298461 639296 298508 639300
rect 298572 639298 298578 639300
rect 298461 639240 298466 639296
rect 298461 639236 298508 639240
rect 298572 639238 298618 639298
rect 298572 639236 298578 639238
rect 298461 639235 298527 639236
rect 301998 638964 302004 639028
rect 302068 639026 302074 639028
rect 373950 639026 374010 639374
rect 381353 639371 381419 639374
rect 381721 639434 381787 639437
rect 385861 639434 385927 639437
rect 381721 639432 385927 639434
rect 381721 639376 381726 639432
rect 381782 639376 385866 639432
rect 385922 639376 385927 639432
rect 381721 639374 385927 639376
rect 381721 639371 381787 639374
rect 385861 639371 385927 639374
rect 302068 638966 374010 639026
rect 302068 638964 302074 638966
rect 49417 637666 49483 637669
rect 49417 637664 52164 637666
rect 49417 637608 49422 637664
rect 49478 637608 52164 637664
rect 49417 637606 52164 637608
rect 49417 637603 49483 637606
rect 478689 636170 478755 636173
rect 478689 636168 480148 636170
rect 478689 636112 478694 636168
rect 478750 636112 480148 636168
rect 478689 636110 480148 636112
rect 478689 636107 478755 636110
rect 254393 634810 254459 634813
rect 251804 634808 254459 634810
rect 251804 634752 254398 634808
rect 254454 634752 254459 634808
rect 251804 634750 254459 634752
rect 254393 634747 254459 634750
rect -960 631940 480 632180
rect 49141 631818 49207 631821
rect 49141 631816 52164 631818
rect 49141 631760 49146 631816
rect 49202 631760 52164 631816
rect 49141 631758 52164 631760
rect 49141 631755 49207 631758
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 521745 630730 521811 630733
rect 519892 630728 521811 630730
rect 519892 630672 521750 630728
rect 521806 630672 521811 630728
rect 583520 630716 584960 630806
rect 519892 630670 521811 630672
rect 521745 630667 521811 630670
rect 278589 630050 278655 630053
rect 278589 630048 280140 630050
rect 278589 629992 278594 630048
rect 278650 629992 280140 630048
rect 278589 629990 280140 629992
rect 278589 629987 278655 629990
rect 254301 628962 254367 628965
rect 251804 628960 254367 628962
rect 251804 628904 254306 628960
rect 254362 628904 254367 628960
rect 251804 628902 254367 628904
rect 254301 628899 254367 628902
rect 50705 625970 50771 625973
rect 50705 625968 52164 625970
rect 50705 625912 50710 625968
rect 50766 625912 52164 625968
rect 50705 625910 52164 625912
rect 50705 625907 50771 625910
rect 254025 623114 254091 623117
rect 251804 623112 254091 623114
rect 251804 623056 254030 623112
rect 254086 623056 254091 623112
rect 251804 623054 254091 623056
rect 254025 623051 254091 623054
rect 48773 620122 48839 620125
rect 48773 620120 52164 620122
rect 48773 620064 48778 620120
rect 48834 620064 52164 620120
rect 48773 620062 52164 620064
rect 48773 620059 48839 620062
rect -960 619170 480 619260
rect -960 619110 674 619170
rect -960 619034 480 619110
rect 614 619034 674 619110
rect -960 619020 674 619034
rect 246 618974 674 619020
rect 246 618490 306 618974
rect 246 618430 6930 618490
rect 6870 618354 6930 618430
rect 50102 618354 50108 618356
rect 6870 618294 50108 618354
rect 50102 618292 50108 618294
rect 50172 618292 50178 618356
rect 478137 617810 478203 617813
rect 478137 617808 480148 617810
rect 478137 617752 478142 617808
rect 478198 617752 480148 617808
rect 478137 617750 480148 617752
rect 478137 617747 478203 617750
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 254669 617266 254735 617269
rect 251804 617264 254735 617266
rect 251804 617208 254674 617264
rect 254730 617208 254735 617264
rect 251804 617206 254735 617208
rect 254669 617203 254735 617206
rect 49182 614212 49188 614276
rect 49252 614274 49258 614276
rect 49252 614214 52164 614274
rect 49252 614212 49258 614214
rect 49182 612716 49188 612780
rect 49252 612778 49258 612780
rect 52085 612778 52151 612781
rect 49252 612776 52151 612778
rect 49252 612720 52090 612776
rect 52146 612720 52151 612776
rect 49252 612718 52151 612720
rect 49252 612716 49258 612718
rect 52085 612715 52151 612718
rect 521653 612370 521719 612373
rect 519892 612368 521719 612370
rect 519892 612312 521658 612368
rect 521714 612312 521719 612368
rect 519892 612310 521719 612312
rect 521653 612307 521719 612310
rect 254485 611418 254551 611421
rect 251804 611416 254551 611418
rect 251804 611360 254490 611416
rect 254546 611360 254551 611416
rect 251804 611358 254551 611360
rect 254485 611355 254551 611358
rect 278681 610058 278747 610061
rect 278681 610056 280140 610058
rect 278681 610000 278686 610056
rect 278742 610000 280140 610056
rect 278681 609998 280140 610000
rect 278681 609995 278747 609998
rect 49366 608364 49372 608428
rect 49436 608426 49442 608428
rect 49436 608366 52164 608426
rect 49436 608364 49442 608366
rect 49366 607140 49372 607204
rect 49436 607202 49442 607204
rect 51993 607202 52059 607205
rect 49436 607200 52059 607202
rect 49436 607144 51998 607200
rect 52054 607144 52059 607200
rect 49436 607142 52059 607144
rect 49436 607140 49442 607142
rect 51993 607139 52059 607142
rect -960 606114 480 606204
rect -960 606054 6930 606114
rect -960 605964 480 606054
rect 6870 605978 6930 606054
rect 49918 605978 49924 605980
rect 6870 605918 49924 605978
rect 49918 605916 49924 605918
rect 49988 605916 49994 605980
rect 254209 605570 254275 605573
rect 251804 605568 254275 605570
rect 251804 605512 254214 605568
rect 254270 605512 254275 605568
rect 251804 605510 254275 605512
rect 254209 605507 254275 605510
rect 583520 604060 584960 604300
rect 49550 602516 49556 602580
rect 49620 602578 49626 602580
rect 49620 602518 52164 602578
rect 49620 602516 49626 602518
rect 49550 600748 49556 600812
rect 49620 600810 49626 600812
rect 51901 600810 51967 600813
rect 49620 600808 51967 600810
rect 49620 600752 51906 600808
rect 51962 600752 51967 600808
rect 49620 600750 51967 600752
rect 49620 600748 49626 600750
rect 51901 600747 51967 600750
rect 301957 600676 302023 600677
rect 303429 600676 303495 600677
rect 301957 600674 302004 600676
rect 301912 600672 302004 600674
rect 301912 600616 301962 600672
rect 301912 600614 302004 600616
rect 301957 600612 302004 600614
rect 302068 600612 302074 600676
rect 303429 600674 303476 600676
rect 303384 600672 303476 600674
rect 303384 600616 303434 600672
rect 303384 600614 303476 600616
rect 303429 600612 303476 600614
rect 303540 600612 303546 600676
rect 306833 600674 306899 600677
rect 307569 600676 307635 600677
rect 307518 600674 307524 600676
rect 306833 600672 307524 600674
rect 307588 600674 307635 600676
rect 307588 600672 307716 600674
rect 306833 600616 306838 600672
rect 306894 600616 307524 600672
rect 307630 600616 307716 600672
rect 306833 600614 307524 600616
rect 301957 600611 302023 600612
rect 303429 600611 303495 600612
rect 306833 600611 306899 600614
rect 307518 600612 307524 600614
rect 307588 600614 307716 600616
rect 307588 600612 307635 600614
rect 307569 600611 307635 600612
rect 254117 599722 254183 599725
rect 251804 599720 254183 599722
rect 251804 599664 254122 599720
rect 254178 599664 254183 599720
rect 251804 599662 254183 599664
rect 254117 599659 254183 599662
rect 302233 598906 302299 598909
rect 302969 598906 303035 598909
rect 302233 598904 303035 598906
rect 302233 598848 302238 598904
rect 302294 598848 302974 598904
rect 303030 598848 303035 598904
rect 302233 598846 303035 598848
rect 302233 598843 302299 598846
rect 302969 598843 303035 598846
rect 360694 598300 360700 598364
rect 360764 598362 360770 598364
rect 370589 598362 370655 598365
rect 360764 598360 370655 598362
rect 360764 598304 370594 598360
rect 370650 598304 370655 598360
rect 360764 598302 370655 598304
rect 360764 598300 360770 598302
rect 370589 598299 370655 598302
rect 300669 598226 300735 598229
rect 319621 598226 319687 598229
rect 300669 598224 319687 598226
rect 300669 598168 300674 598224
rect 300730 598168 319626 598224
rect 319682 598168 319687 598224
rect 300669 598166 319687 598168
rect 300669 598163 300735 598166
rect 319621 598163 319687 598166
rect 366214 598164 366220 598228
rect 366284 598226 366290 598228
rect 367277 598226 367343 598229
rect 366284 598224 367343 598226
rect 366284 598168 367282 598224
rect 367338 598168 367343 598224
rect 366284 598166 367343 598168
rect 366284 598164 366290 598166
rect 367277 598163 367343 598166
rect 369894 598164 369900 598228
rect 369964 598226 369970 598228
rect 371141 598226 371207 598229
rect 369964 598224 371207 598226
rect 369964 598168 371146 598224
rect 371202 598168 371207 598224
rect 369964 598166 371207 598168
rect 369964 598164 369970 598166
rect 371141 598163 371207 598166
rect 378869 598226 378935 598229
rect 379278 598226 379284 598228
rect 378869 598224 379284 598226
rect 378869 598168 378874 598224
rect 378930 598168 379284 598224
rect 378869 598166 379284 598168
rect 378869 598163 378935 598166
rect 379278 598164 379284 598166
rect 379348 598164 379354 598228
rect 373206 597620 373212 597684
rect 373276 597682 373282 597684
rect 376109 597682 376175 597685
rect 373276 597680 376175 597682
rect 373276 597624 376114 597680
rect 376170 597624 376175 597680
rect 373276 597622 376175 597624
rect 373276 597620 373282 597622
rect 376109 597619 376175 597622
rect 362534 596804 362540 596868
rect 362604 596866 362610 596868
rect 391197 596866 391263 596869
rect 362604 596864 391263 596866
rect 362604 596808 391202 596864
rect 391258 596808 391263 596864
rect 362604 596806 391263 596808
rect 362604 596804 362610 596806
rect 391197 596803 391263 596806
rect 404854 596804 404860 596868
rect 404924 596866 404930 596868
rect 479701 596866 479767 596869
rect 404924 596864 479767 596866
rect 404924 596808 479706 596864
rect 479762 596808 479767 596864
rect 404924 596806 479767 596808
rect 404924 596804 404930 596806
rect 479701 596803 479767 596806
rect 48865 596730 48931 596733
rect 48865 596728 52164 596730
rect 48865 596672 48870 596728
rect 48926 596672 52164 596728
rect 48865 596670 52164 596672
rect 48865 596667 48931 596670
rect 382774 595444 382780 595508
rect 382844 595506 382850 595508
rect 392117 595506 392183 595509
rect 382844 595504 392183 595506
rect 382844 595448 392122 595504
rect 392178 595448 392183 595504
rect 382844 595446 392183 595448
rect 382844 595444 382850 595446
rect 392117 595443 392183 595446
rect 254761 593874 254827 593877
rect 251804 593872 254827 593874
rect 251804 593816 254766 593872
rect 254822 593816 254827 593872
rect 251804 593814 254827 593816
rect 254761 593811 254827 593814
rect -960 592908 480 593148
rect 300945 592650 301011 592653
rect 373390 592650 373396 592652
rect 300945 592648 373396 592650
rect 300945 592592 300950 592648
rect 301006 592592 373396 592648
rect 300945 592590 373396 592592
rect 300945 592587 301011 592590
rect 373390 592588 373396 592590
rect 373460 592588 373466 592652
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 48957 590882 49023 590885
rect 48957 590880 52164 590882
rect 48957 590824 48962 590880
rect 49018 590824 52164 590880
rect 583520 590868 584960 590958
rect 48957 590822 52164 590824
rect 48957 590819 49023 590822
rect 254485 588026 254551 588029
rect 251804 588024 254551 588026
rect 251804 587968 254490 588024
rect 254546 587968 254551 588024
rect 251804 587966 254551 587968
rect 254485 587963 254551 587966
rect 395521 586666 395587 586669
rect 394742 586664 395587 586666
rect 394742 586608 395526 586664
rect 395582 586608 395587 586664
rect 394742 586606 395587 586608
rect 392526 586332 392532 586396
rect 392596 586394 392602 586396
rect 394742 586394 394802 586606
rect 395521 586603 395587 586606
rect 392596 586334 394802 586394
rect 392596 586332 392602 586334
rect 364006 585652 364012 585716
rect 364076 585714 364082 585716
rect 396717 585714 396783 585717
rect 364076 585712 396783 585714
rect 364076 585656 396722 585712
rect 396778 585656 396783 585712
rect 364076 585654 396783 585656
rect 364076 585652 364082 585654
rect 396717 585651 396783 585654
rect 48589 585034 48655 585037
rect 48589 585032 52164 585034
rect 48589 584976 48594 585032
rect 48650 584976 52164 585032
rect 48589 584974 52164 584976
rect 48589 584971 48655 584974
rect 387006 583748 387012 583812
rect 387076 583810 387082 583812
rect 389357 583810 389423 583813
rect 387076 583808 389423 583810
rect 387076 583752 389362 583808
rect 389418 583752 389423 583808
rect 387076 583750 389423 583752
rect 387076 583748 387082 583750
rect 389357 583747 389423 583750
rect 362534 583068 362540 583132
rect 362604 583130 362610 583132
rect 378317 583130 378383 583133
rect 362604 583128 378383 583130
rect 362604 583072 378322 583128
rect 378378 583072 378383 583128
rect 362604 583070 378383 583072
rect 362604 583068 362610 583070
rect 378317 583067 378383 583070
rect 299473 582994 299539 582997
rect 388294 582994 388300 582996
rect 299473 582992 388300 582994
rect 299473 582936 299478 582992
rect 299534 582936 388300 582992
rect 299473 582934 388300 582936
rect 299473 582931 299539 582934
rect 388294 582932 388300 582934
rect 388364 582932 388370 582996
rect 253933 582178 253999 582181
rect 251804 582176 253999 582178
rect 251804 582120 253938 582176
rect 253994 582120 253999 582176
rect 251804 582118 253999 582120
rect 253933 582115 253999 582118
rect 379697 581906 379763 581909
rect 391974 581906 391980 581908
rect 379697 581904 391980 581906
rect 379697 581848 379702 581904
rect 379758 581848 391980 581904
rect 379697 581846 391980 581848
rect 379697 581843 379763 581846
rect 391974 581844 391980 581846
rect 392044 581844 392050 581908
rect 368238 581708 368244 581772
rect 368308 581770 368314 581772
rect 382457 581770 382523 581773
rect 368308 581768 382523 581770
rect 368308 581712 382462 581768
rect 382518 581712 382523 581768
rect 368308 581710 382523 581712
rect 368308 581708 368314 581710
rect 382457 581707 382523 581710
rect 300669 581634 300735 581637
rect 380934 581634 380940 581636
rect 300669 581632 380940 581634
rect 300669 581576 300674 581632
rect 300730 581576 380940 581632
rect 300669 581574 380940 581576
rect 300669 581571 300735 581574
rect 380934 581572 380940 581574
rect 381004 581572 381010 581636
rect 371734 580348 371740 580412
rect 371804 580410 371810 580412
rect 386597 580410 386663 580413
rect 371804 580408 386663 580410
rect 371804 580352 386602 580408
rect 386658 580352 386663 580408
rect 371804 580350 386663 580352
rect 371804 580348 371810 580350
rect 386597 580347 386663 580350
rect 299381 580274 299447 580277
rect 376150 580274 376156 580276
rect 299381 580272 376156 580274
rect 299381 580216 299386 580272
rect 299442 580216 376156 580272
rect 299381 580214 376156 580216
rect 299381 580211 299447 580214
rect 376150 580212 376156 580214
rect 376220 580212 376226 580276
rect -960 579852 480 580092
rect 48681 579186 48747 579189
rect 48681 579184 52164 579186
rect 48681 579128 48686 579184
rect 48742 579128 52164 579184
rect 48681 579126 52164 579128
rect 48681 579123 48747 579126
rect 282678 578988 282684 579052
rect 282748 579050 282754 579052
rect 473997 579050 474063 579053
rect 282748 579048 474063 579050
rect 282748 578992 474002 579048
rect 474058 578992 474063 579048
rect 282748 578990 474063 578992
rect 282748 578988 282754 578990
rect 473997 578987 474063 578990
rect 311014 578852 311020 578916
rect 311084 578914 311090 578916
rect 580257 578914 580323 578917
rect 311084 578912 580323 578914
rect 311084 578856 580262 578912
rect 580318 578856 580323 578912
rect 311084 578854 580323 578856
rect 311084 578852 311090 578854
rect 580257 578851 580323 578854
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 376753 576874 376819 576877
rect 384062 576874 384068 576876
rect 376753 576872 384068 576874
rect 376753 576816 376758 576872
rect 376814 576816 384068 576872
rect 376753 576814 384068 576816
rect 376753 576811 376819 576814
rect 384062 576812 384068 576814
rect 384132 576812 384138 576876
rect 254485 576330 254551 576333
rect 251804 576328 254551 576330
rect 251804 576272 254490 576328
rect 254546 576272 254551 576328
rect 251804 576270 254551 576272
rect 254485 576267 254551 576270
rect 292665 574834 292731 574837
rect 391054 574834 391060 574836
rect 292665 574832 391060 574834
rect 292665 574776 292670 574832
rect 292726 574776 391060 574832
rect 292665 574774 391060 574776
rect 292665 574771 292731 574774
rect 391054 574772 391060 574774
rect 391124 574772 391130 574836
rect 287053 574698 287119 574701
rect 389582 574698 389588 574700
rect 287053 574696 389588 574698
rect 287053 574640 287058 574696
rect 287114 574640 389588 574696
rect 287053 574638 389588 574640
rect 287053 574635 287119 574638
rect 389582 574636 389588 574638
rect 389652 574636 389658 574700
rect 49325 573338 49391 573341
rect 281625 573338 281691 573341
rect 396574 573338 396580 573340
rect 49325 573336 52164 573338
rect 49325 573280 49330 573336
rect 49386 573280 52164 573336
rect 49325 573278 52164 573280
rect 281625 573336 396580 573338
rect 281625 573280 281630 573336
rect 281686 573280 396580 573336
rect 281625 573278 396580 573280
rect 49325 573275 49391 573278
rect 281625 573275 281691 573278
rect 396574 573276 396580 573278
rect 396644 573276 396650 573340
rect 284293 571978 284359 571981
rect 370078 571978 370084 571980
rect 284293 571976 370084 571978
rect 284293 571920 284298 571976
rect 284354 571920 370084 571976
rect 284293 571918 370084 571920
rect 284293 571915 284359 571918
rect 370078 571916 370084 571918
rect 370148 571916 370154 571980
rect 253933 570482 253999 570485
rect 251804 570480 253999 570482
rect 251804 570424 253938 570480
rect 253994 570424 253999 570480
rect 251804 570422 253999 570424
rect 253933 570419 253999 570422
rect 362350 569196 362356 569260
rect 362420 569258 362426 569260
rect 369945 569258 370011 569261
rect 362420 569256 370011 569258
rect 362420 569200 369950 569256
rect 370006 569200 370011 569256
rect 362420 569198 370011 569200
rect 362420 569196 362426 569198
rect 369945 569195 370011 569198
rect 311893 568170 311959 568173
rect 376886 568170 376892 568172
rect 311893 568168 376892 568170
rect 311893 568112 311898 568168
rect 311954 568112 376892 568168
rect 311893 568110 376892 568112
rect 311893 568107 311959 568110
rect 376886 568108 376892 568110
rect 376956 568108 376962 568172
rect 294597 568034 294663 568037
rect 368422 568034 368428 568036
rect 294597 568032 368428 568034
rect 294597 567976 294602 568032
rect 294658 567976 368428 568032
rect 294597 567974 368428 567976
rect 294597 567971 294663 567974
rect 368422 567972 368428 567974
rect 368492 567972 368498 568036
rect 376334 567972 376340 568036
rect 376404 568034 376410 568036
rect 388529 568034 388595 568037
rect 376404 568032 388595 568034
rect 376404 567976 388534 568032
rect 388590 567976 388595 568032
rect 376404 567974 388595 567976
rect 376404 567972 376410 567974
rect 388529 567971 388595 567974
rect 279366 567836 279372 567900
rect 279436 567898 279442 567900
rect 512177 567898 512243 567901
rect 279436 567896 512243 567898
rect 279436 567840 512182 567896
rect 512238 567840 512243 567896
rect 279436 567838 512243 567840
rect 279436 567836 279442 567838
rect 512177 567835 512243 567838
rect 49049 567490 49115 567493
rect 49049 567488 52164 567490
rect 49049 567432 49054 567488
rect 49110 567432 52164 567488
rect 49049 567430 52164 567432
rect 49049 567427 49115 567430
rect -960 566946 480 567036
rect -960 566886 674 566946
rect -960 566810 480 566886
rect 614 566810 674 566886
rect -960 566796 674 566810
rect 246 566750 674 566796
rect 246 566266 306 566750
rect 319437 566402 319503 566405
rect 380566 566402 380572 566404
rect 319437 566400 380572 566402
rect 319437 566344 319442 566400
rect 319498 566344 380572 566400
rect 319437 566342 380572 566344
rect 319437 566339 319503 566342
rect 380566 566340 380572 566342
rect 380636 566340 380642 566404
rect 246 566206 6930 566266
rect 6870 565858 6930 566206
rect 49734 565858 49740 565860
rect 6870 565798 49740 565858
rect 49734 565796 49740 565798
rect 49804 565796 49810 565860
rect 361614 565116 361620 565180
rect 361684 565178 361690 565180
rect 382365 565178 382431 565181
rect 361684 565176 382431 565178
rect 361684 565120 382370 565176
rect 382426 565120 382431 565176
rect 361684 565118 382431 565120
rect 361684 565116 361690 565118
rect 382365 565115 382431 565118
rect 320909 565042 320975 565045
rect 373758 565042 373764 565044
rect 320909 565040 373764 565042
rect 320909 564984 320914 565040
rect 320970 564984 373764 565040
rect 320909 564982 373764 564984
rect 320909 564979 320975 564982
rect 373758 564980 373764 564982
rect 373828 564980 373834 565044
rect 279366 564634 279372 564636
rect 251804 564574 279372 564634
rect 279366 564572 279372 564574
rect 279436 564572 279442 564636
rect 580349 564362 580415 564365
rect 583520 564362 584960 564452
rect 580349 564360 584960 564362
rect 580349 564304 580354 564360
rect 580410 564304 584960 564360
rect 580349 564302 584960 564304
rect 580349 564299 580415 564302
rect 583520 564212 584960 564302
rect 361430 563892 361436 563956
rect 361500 563954 361506 563956
rect 378225 563954 378291 563957
rect 361500 563952 378291 563954
rect 361500 563896 378230 563952
rect 378286 563896 378291 563952
rect 361500 563894 378291 563896
rect 361500 563892 361506 563894
rect 378225 563891 378291 563894
rect 309317 563818 309383 563821
rect 400254 563818 400260 563820
rect 309317 563816 400260 563818
rect 309317 563760 309322 563816
rect 309378 563760 400260 563816
rect 309317 563758 400260 563760
rect 309317 563755 309383 563758
rect 400254 563756 400260 563758
rect 400324 563756 400330 563820
rect 285438 563620 285444 563684
rect 285508 563682 285514 563684
rect 398782 563682 398788 563684
rect 285508 563622 398788 563682
rect 285508 563620 285514 563622
rect 398782 563620 398788 563622
rect 398852 563620 398858 563684
rect 298318 562260 298324 562324
rect 298388 562322 298394 562324
rect 399150 562322 399156 562324
rect 298388 562262 399156 562322
rect 298388 562260 298394 562262
rect 399150 562260 399156 562262
rect 399220 562260 399226 562324
rect 49233 561642 49299 561645
rect 49233 561640 52164 561642
rect 49233 561584 49238 561640
rect 49294 561584 52164 561640
rect 49233 561582 52164 561584
rect 49233 561579 49299 561582
rect 362718 561036 362724 561100
rect 362788 561098 362794 561100
rect 400489 561098 400555 561101
rect 362788 561096 400555 561098
rect 362788 561040 400494 561096
rect 400550 561040 400555 561096
rect 362788 561038 400555 561040
rect 362788 561036 362794 561038
rect 400489 561035 400555 561038
rect 282913 560962 282979 560965
rect 364742 560962 364748 560964
rect 282913 560960 364748 560962
rect 282913 560904 282918 560960
rect 282974 560904 364748 560960
rect 282913 560902 364748 560904
rect 282913 560899 282979 560902
rect 364742 560900 364748 560902
rect 364812 560900 364818 560964
rect 361665 560282 361731 560285
rect 362902 560282 362908 560284
rect 361665 560280 362908 560282
rect 361665 560224 361670 560280
rect 361726 560224 362908 560280
rect 361665 560222 362908 560224
rect 361665 560219 361731 560222
rect 362902 560220 362908 560222
rect 362972 560220 362978 560284
rect 385534 560220 385540 560284
rect 385604 560282 385610 560284
rect 388437 560282 388503 560285
rect 385604 560280 388503 560282
rect 385604 560224 388442 560280
rect 388498 560224 388503 560280
rect 385604 560222 388503 560224
rect 385604 560220 385610 560222
rect 388437 560219 388503 560222
rect 298502 559540 298508 559604
rect 298572 559602 298578 559604
rect 399569 559602 399635 559605
rect 298572 559600 399635 559602
rect 298572 559544 399574 559600
rect 399630 559544 399635 559600
rect 298572 559542 399635 559544
rect 298572 559540 298578 559542
rect 399569 559539 399635 559542
rect 361757 558922 361823 558925
rect 363454 558922 363460 558924
rect 361757 558920 363460 558922
rect 361757 558864 361762 558920
rect 361818 558864 363460 558920
rect 361757 558862 363460 558864
rect 361757 558859 361823 558862
rect 363454 558860 363460 558862
rect 363524 558860 363530 558924
rect 254577 558786 254643 558789
rect 251804 558784 254643 558786
rect 251804 558728 254582 558784
rect 254638 558728 254643 558784
rect 251804 558726 254643 558728
rect 254577 558723 254643 558726
rect 314653 558242 314719 558245
rect 400438 558242 400444 558244
rect 314653 558240 400444 558242
rect 314653 558184 314658 558240
rect 314714 558184 400444 558240
rect 314653 558182 400444 558184
rect 314653 558179 314719 558182
rect 400438 558180 400444 558182
rect 400508 558180 400514 558244
rect 48773 555794 48839 555797
rect 48773 555792 52164 555794
rect 48773 555736 48778 555792
rect 48834 555736 52164 555792
rect 48773 555734 52164 555736
rect 48773 555731 48839 555734
rect 321001 555386 321067 555389
rect 401726 555386 401732 555388
rect 321001 555384 401732 555386
rect 321001 555328 321006 555384
rect 321062 555328 401732 555384
rect 321001 555326 401732 555328
rect 321001 555323 321067 555326
rect 401726 555324 401732 555326
rect 401796 555324 401802 555388
rect 359038 554236 359044 554300
rect 359108 554298 359114 554300
rect 368473 554298 368539 554301
rect 359108 554296 368539 554298
rect 359108 554240 368478 554296
rect 368534 554240 368539 554296
rect 359108 554238 368539 554240
rect 359108 554236 359114 554238
rect 368473 554235 368539 554238
rect 289486 554100 289492 554164
rect 289556 554162 289562 554164
rect 400622 554162 400628 554164
rect 289556 554102 400628 554162
rect 289556 554100 289562 554102
rect 400622 554100 400628 554102
rect 400692 554100 400698 554164
rect -960 553890 480 553980
rect 358854 553964 358860 554028
rect 358924 554026 358930 554028
rect 580349 554026 580415 554029
rect 358924 554024 580415 554026
rect 358924 553968 580354 554024
rect 580410 553968 580415 554024
rect 358924 553966 580415 553968
rect 358924 553964 358930 553966
rect 580349 553963 580415 553966
rect 3785 553890 3851 553893
rect -960 553888 3851 553890
rect -960 553832 3790 553888
rect 3846 553832 3851 553888
rect -960 553830 3851 553832
rect -960 553740 480 553830
rect 3785 553827 3851 553830
rect 358302 553420 358308 553484
rect 358372 553482 358378 553484
rect 363597 553482 363663 553485
rect 358372 553480 363663 553482
rect 358372 553424 363602 553480
rect 363658 553424 363663 553480
rect 358372 553422 363663 553424
rect 358372 553420 358378 553422
rect 363597 553419 363663 553422
rect 254393 552938 254459 552941
rect 251804 552936 254459 552938
rect 251804 552880 254398 552936
rect 254454 552880 254459 552936
rect 251804 552878 254459 552880
rect 254393 552875 254459 552878
rect 369025 552122 369091 552125
rect 403566 552122 403572 552124
rect 369025 552120 403572 552122
rect 369025 552064 369030 552120
rect 369086 552064 403572 552120
rect 369025 552062 403572 552064
rect 369025 552059 369091 552062
rect 403566 552060 403572 552062
rect 403636 552060 403642 552124
rect 358670 551924 358676 551988
rect 358740 551986 358746 551988
rect 360929 551986 360995 551989
rect 358740 551984 360995 551986
rect 358740 551928 360934 551984
rect 360990 551928 360995 551984
rect 358740 551926 360995 551928
rect 358740 551924 358746 551926
rect 360929 551923 360995 551926
rect 358486 551788 358492 551852
rect 358556 551850 358562 551852
rect 361573 551850 361639 551853
rect 358556 551848 361639 551850
rect 358556 551792 361578 551848
rect 361634 551792 361639 551848
rect 358556 551790 361639 551792
rect 358556 551788 358562 551790
rect 361573 551787 361639 551790
rect 293166 551516 293172 551580
rect 293236 551578 293242 551580
rect 401685 551578 401751 551581
rect 293236 551576 401751 551578
rect 293236 551520 401690 551576
rect 401746 551520 401751 551576
rect 293236 551518 401751 551520
rect 293236 551516 293242 551518
rect 401685 551515 401751 551518
rect 288198 551380 288204 551444
rect 288268 551442 288274 551444
rect 400806 551442 400812 551444
rect 288268 551382 400812 551442
rect 288268 551380 288274 551382
rect 400806 551380 400812 551382
rect 400876 551380 400882 551444
rect 280153 551306 280219 551309
rect 398966 551306 398972 551308
rect 280153 551304 398972 551306
rect 280153 551248 280158 551304
rect 280214 551248 398972 551304
rect 280153 551246 398972 551248
rect 280153 551243 280219 551246
rect 398966 551244 398972 551246
rect 399036 551244 399042 551308
rect 583520 551020 584960 551260
rect 358118 550564 358124 550628
rect 358188 550626 358194 550628
rect 360837 550626 360903 550629
rect 358188 550624 360903 550626
rect 358188 550568 360842 550624
rect 360898 550568 360903 550624
rect 358188 550566 360903 550568
rect 358188 550564 358194 550566
rect 360837 550563 360903 550566
rect 397453 550626 397519 550629
rect 398097 550626 398163 550629
rect 399334 550626 399340 550628
rect 397453 550624 399340 550626
rect 397453 550568 397458 550624
rect 397514 550568 398102 550624
rect 398158 550568 399340 550624
rect 397453 550566 399340 550568
rect 397453 550563 397519 550566
rect 398097 550563 398163 550566
rect 399334 550564 399340 550566
rect 399404 550564 399410 550628
rect 357157 550354 357223 550357
rect 357157 550352 360210 550354
rect 357157 550296 357162 550352
rect 357218 550296 360210 550352
rect 357157 550294 360210 550296
rect 357157 550291 357223 550294
rect 49141 549946 49207 549949
rect 49141 549944 52164 549946
rect 49141 549888 49146 549944
rect 49202 549888 52164 549944
rect 49141 549886 52164 549888
rect 49141 549883 49207 549886
rect 360150 549712 360210 550294
rect 401542 549266 401548 549268
rect 399894 549206 401548 549266
rect 399894 549032 399954 549206
rect 401542 549204 401548 549206
rect 401612 549204 401618 549268
rect 357617 548586 357683 548589
rect 360150 548586 360210 549032
rect 357617 548584 360210 548586
rect 357617 548528 357622 548584
rect 357678 548528 360210 548584
rect 357617 548526 360210 548528
rect 357617 548523 357683 548526
rect 357893 548450 357959 548453
rect 357893 548448 360210 548450
rect 357893 548392 357898 548448
rect 357954 548392 360210 548448
rect 357893 548390 360210 548392
rect 357893 548387 357959 548390
rect 360150 548352 360210 548390
rect 357433 547770 357499 547773
rect 400806 547770 400812 547772
rect 357433 547768 360210 547770
rect 357433 547712 357438 547768
rect 357494 547712 360210 547768
rect 357433 547710 360210 547712
rect 357433 547707 357499 547710
rect 360150 547672 360210 547710
rect 399894 547710 400812 547770
rect 399894 547672 399954 547710
rect 400806 547708 400812 547710
rect 400876 547708 400882 547772
rect 401593 547498 401659 547501
rect 399894 547496 401659 547498
rect 399894 547440 401598 547496
rect 401654 547440 401659 547496
rect 399894 547438 401659 547440
rect 254485 547090 254551 547093
rect 251804 547088 254551 547090
rect 251804 547032 254490 547088
rect 254546 547032 254551 547088
rect 251804 547030 254551 547032
rect 254485 547027 254551 547030
rect 332041 547090 332107 547093
rect 358302 547090 358308 547092
rect 332041 547088 358308 547090
rect 332041 547032 332046 547088
rect 332102 547032 358308 547088
rect 332041 547030 358308 547032
rect 332041 547027 332107 547030
rect 358302 547028 358308 547030
rect 358372 547090 358378 547092
rect 358372 547030 360210 547090
rect 358372 547028 358378 547030
rect 360150 546992 360210 547030
rect 399894 546992 399954 547438
rect 401593 547435 401659 547438
rect 403065 546410 403131 546413
rect 399894 546408 403131 546410
rect 399894 546352 403070 546408
rect 403126 546352 403131 546408
rect 399894 546350 403131 546352
rect 399894 546312 399954 546350
rect 403065 546347 403131 546350
rect 399937 546138 400003 546141
rect 399894 546136 400003 546138
rect 399894 546080 399942 546136
rect 399998 546080 400003 546136
rect 399894 546075 400003 546080
rect 357433 546002 357499 546005
rect 357433 546000 360210 546002
rect 357433 545944 357438 546000
rect 357494 545944 360210 546000
rect 357433 545942 360210 545944
rect 357433 545939 357499 545942
rect 360150 545632 360210 545942
rect 399894 545632 399954 546075
rect 358721 545050 358787 545053
rect 358721 545048 360210 545050
rect 358721 544992 358726 545048
rect 358782 544992 360210 545048
rect 358721 544990 360210 544992
rect 358721 544987 358787 544990
rect 360150 544952 360210 544990
rect 401685 544778 401751 544781
rect 399894 544776 401751 544778
rect 399894 544720 401690 544776
rect 401746 544720 401751 544776
rect 399894 544718 401751 544720
rect 357433 544642 357499 544645
rect 357433 544640 360210 544642
rect 357433 544584 357438 544640
rect 357494 544584 360210 544640
rect 357433 544582 360210 544584
rect 357433 544579 357499 544582
rect 360150 544272 360210 544582
rect 399894 544272 399954 544718
rect 401685 544715 401751 544718
rect 49417 544098 49483 544101
rect 49417 544096 52164 544098
rect 49417 544040 49422 544096
rect 49478 544040 52164 544096
rect 49417 544038 52164 544040
rect 49417 544035 49483 544038
rect 399334 543764 399340 543828
rect 399404 543764 399410 543828
rect 317505 543690 317571 543693
rect 317638 543690 317644 543692
rect 317505 543688 317644 543690
rect 317505 543632 317510 543688
rect 317566 543632 317644 543688
rect 317505 543630 317644 543632
rect 317505 543627 317571 543630
rect 317638 543628 317644 543630
rect 317708 543628 317714 543692
rect 399342 543592 399402 543764
rect 357525 543554 357591 543557
rect 357985 543554 358051 543557
rect 360150 543554 360210 543592
rect 357525 543552 360210 543554
rect 357525 543496 357530 543552
rect 357586 543496 357990 543552
rect 358046 543496 360210 543552
rect 357525 543494 360210 543496
rect 357525 543491 357591 543494
rect 357985 543491 358051 543494
rect 290958 543356 290964 543420
rect 291028 543418 291034 543420
rect 296161 543418 296227 543421
rect 291028 543416 296227 543418
rect 291028 543360 296166 543416
rect 296222 543360 296227 543416
rect 291028 543358 296227 543360
rect 291028 543356 291034 543358
rect 296161 543355 296227 543358
rect 358813 543418 358879 543421
rect 358813 543416 360210 543418
rect 358813 543360 358818 543416
rect 358874 543360 360210 543416
rect 358813 543358 360210 543360
rect 358813 543355 358879 543358
rect 295926 543220 295932 543284
rect 295996 543282 296002 543284
rect 307017 543282 307083 543285
rect 295996 543280 307083 543282
rect 295996 543224 307022 543280
rect 307078 543224 307083 543280
rect 295996 543222 307083 543224
rect 295996 543220 296002 543222
rect 307017 543219 307083 543222
rect 286174 543084 286180 543148
rect 286244 543146 286250 543148
rect 301865 543146 301931 543149
rect 286244 543144 301931 543146
rect 286244 543088 301870 543144
rect 301926 543088 301931 543144
rect 286244 543086 301931 543088
rect 286244 543084 286250 543086
rect 301865 543083 301931 543086
rect 283414 542948 283420 543012
rect 283484 543010 283490 543012
rect 283484 542950 302250 543010
rect 283484 542948 283490 542950
rect 291694 542812 291700 542876
rect 291764 542874 291770 542876
rect 298185 542874 298251 542877
rect 291764 542872 298251 542874
rect 291764 542816 298190 542872
rect 298246 542816 298251 542872
rect 291764 542814 298251 542816
rect 302190 542874 302250 542950
rect 360150 542912 360210 543358
rect 401593 543146 401659 543149
rect 399894 543144 401659 543146
rect 399894 543088 401598 543144
rect 401654 543088 401659 543144
rect 399894 543086 401659 543088
rect 399894 542912 399954 543086
rect 401593 543083 401659 543086
rect 304073 542874 304139 542877
rect 302190 542872 304139 542874
rect 302190 542816 304078 542872
rect 304134 542816 304139 542872
rect 302190 542814 304139 542816
rect 291764 542812 291770 542814
rect 298185 542811 298251 542814
rect 304073 542811 304139 542814
rect 311934 542812 311940 542876
rect 312004 542874 312010 542876
rect 312261 542874 312327 542877
rect 312004 542872 312327 542874
rect 312004 542816 312266 542872
rect 312322 542816 312327 542872
rect 312004 542814 312327 542816
rect 312004 542812 312010 542814
rect 312261 542811 312327 542814
rect 279785 542738 279851 542741
rect 292573 542738 292639 542741
rect 279785 542736 292639 542738
rect 279785 542680 279790 542736
rect 279846 542680 292578 542736
rect 292634 542680 292639 542736
rect 279785 542678 292639 542680
rect 279785 542675 279851 542678
rect 292573 542675 292639 542678
rect 296161 542738 296227 542741
rect 304993 542738 305059 542741
rect 296161 542736 305059 542738
rect 296161 542680 296166 542736
rect 296222 542680 304998 542736
rect 305054 542680 305059 542736
rect 296161 542678 305059 542680
rect 296161 542675 296227 542678
rect 304993 542675 305059 542678
rect 308622 542676 308628 542740
rect 308692 542738 308698 542740
rect 310697 542738 310763 542741
rect 308692 542736 310763 542738
rect 308692 542680 310702 542736
rect 310758 542680 310763 542736
rect 308692 542678 310763 542680
rect 308692 542676 308698 542678
rect 310697 542675 310763 542678
rect 295006 542540 295012 542604
rect 295076 542602 295082 542604
rect 298921 542602 298987 542605
rect 295076 542600 298987 542602
rect 295076 542544 298926 542600
rect 298982 542544 298987 542600
rect 295076 542542 298987 542544
rect 295076 542540 295082 542542
rect 298921 542539 298987 542542
rect 305494 542540 305500 542604
rect 305564 542602 305570 542604
rect 308489 542602 308555 542605
rect 305564 542600 308555 542602
rect 305564 542544 308494 542600
rect 308550 542544 308555 542600
rect 305564 542542 308555 542544
rect 305564 542540 305570 542542
rect 308489 542539 308555 542542
rect 309358 542540 309364 542604
rect 309428 542602 309434 542604
rect 309961 542602 310027 542605
rect 309428 542600 310027 542602
rect 309428 542544 309966 542600
rect 310022 542544 310027 542600
rect 309428 542542 310027 542544
rect 309428 542540 309434 542542
rect 309961 542539 310027 542542
rect 297173 542468 297239 542469
rect 299933 542468 299999 542469
rect 297173 542466 297220 542468
rect 297128 542464 297220 542466
rect 297128 542408 297178 542464
rect 297128 542406 297220 542408
rect 297173 542404 297220 542406
rect 297284 542404 297290 542468
rect 299933 542466 299980 542468
rect 299888 542464 299980 542466
rect 299888 542408 299938 542464
rect 299888 542406 299980 542408
rect 299933 542404 299980 542406
rect 300044 542404 300050 542468
rect 304206 542404 304212 542468
rect 304276 542466 304282 542468
rect 306373 542466 306439 542469
rect 304276 542464 306439 542466
rect 304276 542408 306378 542464
rect 306434 542408 306439 542464
rect 304276 542406 306439 542408
rect 304276 542404 304282 542406
rect 297173 542403 297239 542404
rect 299933 542403 299999 542404
rect 306373 542403 306439 542406
rect 308397 542466 308463 542469
rect 308806 542466 308812 542468
rect 308397 542464 308812 542466
rect 308397 542408 308402 542464
rect 308458 542408 308812 542464
rect 308397 542406 308812 542408
rect 308397 542403 308463 542406
rect 308806 542404 308812 542406
rect 308876 542404 308882 542468
rect 309174 542404 309180 542468
rect 309244 542466 309250 542468
rect 309409 542466 309475 542469
rect 309244 542464 309475 542466
rect 309244 542408 309414 542464
rect 309470 542408 309475 542464
rect 309244 542406 309475 542408
rect 309244 542404 309250 542406
rect 309409 542403 309475 542406
rect 310462 542404 310468 542468
rect 310532 542466 310538 542468
rect 311433 542466 311499 542469
rect 310532 542464 311499 542466
rect 310532 542408 311438 542464
rect 311494 542408 311499 542464
rect 310532 542406 311499 542408
rect 310532 542404 310538 542406
rect 311433 542403 311499 542406
rect 359181 542330 359247 542333
rect 359181 542328 360210 542330
rect 359181 542272 359186 542328
rect 359242 542272 360210 542328
rect 359181 542270 360210 542272
rect 359181 542267 359247 542270
rect 360150 542232 360210 542270
rect 399894 541786 399954 542232
rect 401593 541786 401659 541789
rect 399894 541784 401659 541786
rect 399894 541728 401598 541784
rect 401654 541728 401659 541784
rect 399894 541726 401659 541728
rect 401593 541723 401659 541726
rect 400121 541582 400187 541585
rect 399924 541580 400187 541582
rect 254577 541242 254643 541245
rect 251804 541240 254643 541242
rect 251804 541184 254582 541240
rect 254638 541184 254643 541240
rect 251804 541182 254643 541184
rect 254577 541179 254643 541182
rect 327901 541106 327967 541109
rect 359038 541106 359044 541108
rect 327901 541104 359044 541106
rect 327901 541048 327906 541104
rect 327962 541048 359044 541104
rect 327901 541046 359044 541048
rect 327901 541043 327967 541046
rect 359038 541044 359044 541046
rect 359108 541106 359114 541108
rect 360150 541106 360210 541552
rect 399924 541524 400126 541580
rect 400182 541524 400187 541580
rect 399924 541522 400187 541524
rect 400121 541519 400187 541522
rect 359108 541046 360210 541106
rect 359108 541044 359114 541046
rect 358445 540970 358511 540973
rect 401961 540970 402027 540973
rect 358445 540968 360210 540970
rect -960 540684 480 540924
rect 358445 540912 358450 540968
rect 358506 540912 360210 540968
rect 358445 540910 360210 540912
rect 358445 540907 358511 540910
rect 360150 540872 360210 540910
rect 399894 540968 402027 540970
rect 399894 540912 401966 540968
rect 402022 540912 402027 540968
rect 399894 540910 402027 540912
rect 399894 540872 399954 540910
rect 401961 540907 402027 540910
rect 358118 540636 358124 540700
rect 358188 540698 358194 540700
rect 400949 540698 401015 540701
rect 358188 540638 360210 540698
rect 358188 540636 358194 540638
rect 360150 540192 360210 540638
rect 399894 540696 401015 540698
rect 399894 540640 400954 540696
rect 401010 540640 401015 540696
rect 399894 540638 401015 540640
rect 399894 540192 399954 540638
rect 400949 540635 401015 540638
rect 287278 539684 287284 539748
rect 287348 539746 287354 539748
rect 287881 539746 287947 539749
rect 287348 539744 287947 539746
rect 287348 539688 287886 539744
rect 287942 539688 287947 539744
rect 287348 539686 287947 539688
rect 287348 539684 287354 539686
rect 287881 539683 287947 539686
rect 49182 539548 49188 539612
rect 49252 539610 49258 539612
rect 49417 539610 49483 539613
rect 49252 539608 49483 539610
rect 49252 539552 49422 539608
rect 49478 539552 49483 539608
rect 49252 539550 49483 539552
rect 49252 539548 49258 539550
rect 49417 539547 49483 539550
rect 283373 539610 283439 539613
rect 284886 539610 284892 539612
rect 283373 539608 284892 539610
rect 283373 539552 283378 539608
rect 283434 539552 284892 539608
rect 283373 539550 284892 539552
rect 283373 539547 283439 539550
rect 284886 539548 284892 539550
rect 284956 539548 284962 539612
rect 285990 539548 285996 539612
rect 286060 539610 286066 539612
rect 286133 539610 286199 539613
rect 286060 539608 286199 539610
rect 286060 539552 286138 539608
rect 286194 539552 286199 539608
rect 286060 539550 286199 539552
rect 286060 539548 286066 539550
rect 286133 539547 286199 539550
rect 287462 539548 287468 539612
rect 287532 539610 287538 539612
rect 287605 539610 287671 539613
rect 287532 539608 287671 539610
rect 287532 539552 287610 539608
rect 287666 539552 287671 539608
rect 287532 539550 287671 539552
rect 287532 539548 287538 539550
rect 287605 539547 287671 539550
rect 288382 539548 288388 539612
rect 288452 539610 288458 539612
rect 288617 539610 288683 539613
rect 288452 539608 288683 539610
rect 288452 539552 288622 539608
rect 288678 539552 288683 539608
rect 288452 539550 288683 539552
rect 288452 539548 288458 539550
rect 288617 539547 288683 539550
rect 288750 539548 288756 539612
rect 288820 539610 288826 539612
rect 289353 539610 289419 539613
rect 288820 539608 289419 539610
rect 288820 539552 289358 539608
rect 289414 539552 289419 539608
rect 288820 539550 289419 539552
rect 288820 539548 288826 539550
rect 289353 539547 289419 539550
rect 290549 539612 290615 539613
rect 290825 539612 290891 539613
rect 290549 539608 290596 539612
rect 290660 539610 290666 539612
rect 290549 539552 290554 539608
rect 290549 539548 290596 539552
rect 290660 539550 290706 539610
rect 290660 539548 290666 539550
rect 290774 539548 290780 539612
rect 290844 539610 290891 539612
rect 290844 539608 290936 539610
rect 290886 539552 290936 539608
rect 290844 539550 290936 539552
rect 290844 539548 290891 539550
rect 291142 539548 291148 539612
rect 291212 539610 291218 539612
rect 291561 539610 291627 539613
rect 291212 539608 291627 539610
rect 291212 539552 291566 539608
rect 291622 539552 291627 539608
rect 291212 539550 291627 539552
rect 291212 539548 291218 539550
rect 290549 539547 290615 539548
rect 290825 539547 290891 539548
rect 291561 539547 291627 539550
rect 292798 539548 292804 539612
rect 292868 539610 292874 539612
rect 293033 539610 293099 539613
rect 403014 539610 403020 539612
rect 292868 539608 293099 539610
rect 292868 539552 293038 539608
rect 293094 539552 293099 539608
rect 292868 539550 293099 539552
rect 292868 539548 292874 539550
rect 293033 539547 293099 539550
rect 399894 539550 403020 539610
rect 399894 539512 399954 539550
rect 403014 539548 403020 539550
rect 403084 539548 403090 539612
rect 358813 539338 358879 539341
rect 360150 539338 360210 539512
rect 401041 539338 401107 539341
rect 358813 539336 360210 539338
rect 358813 539280 358818 539336
rect 358874 539280 360210 539336
rect 358813 539278 360210 539280
rect 399894 539336 401107 539338
rect 399894 539280 401046 539336
rect 401102 539280 401107 539336
rect 399894 539278 401107 539280
rect 358813 539275 358879 539278
rect 357433 539202 357499 539205
rect 357433 539200 360210 539202
rect 357433 539144 357438 539200
rect 357494 539144 360210 539200
rect 357433 539142 360210 539144
rect 357433 539139 357499 539142
rect 360150 538832 360210 539142
rect 399894 538832 399954 539278
rect 401041 539275 401107 539278
rect 49417 538250 49483 538253
rect 49417 538248 52164 538250
rect 49417 538192 49422 538248
rect 49478 538192 52164 538248
rect 49417 538190 52164 538192
rect 49417 538187 49483 538190
rect 358353 538114 358419 538117
rect 360150 538114 360210 538152
rect 358353 538112 360210 538114
rect 358353 538056 358358 538112
rect 358414 538056 360210 538112
rect 358353 538054 360210 538056
rect 399894 538114 399954 538152
rect 400765 538114 400831 538117
rect 399894 538112 400831 538114
rect 399894 538056 400770 538112
rect 400826 538056 400831 538112
rect 399894 538054 400831 538056
rect 358353 538051 358419 538054
rect 400765 538051 400831 538054
rect 358905 537842 358971 537845
rect 400622 537842 400628 537844
rect 358905 537840 360210 537842
rect 358905 537784 358910 537840
rect 358966 537784 360210 537840
rect 358905 537782 360210 537784
rect 358905 537779 358971 537782
rect 360150 537472 360210 537782
rect 399894 537782 400628 537842
rect 399894 537472 399954 537782
rect 400622 537780 400628 537782
rect 400692 537780 400698 537844
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect 320173 537366 320239 537369
rect 319884 537364 320239 537366
rect 319884 537308 320178 537364
rect 320234 537308 320239 537364
rect 319884 537306 320239 537308
rect 320173 537303 320239 537306
rect 357433 536754 357499 536757
rect 360150 536754 360210 536792
rect 357433 536752 360210 536754
rect 357433 536696 357438 536752
rect 357494 536696 360210 536752
rect 357433 536694 360210 536696
rect 357433 536691 357499 536694
rect 319854 536210 319914 536656
rect 399894 536621 399954 536792
rect 357893 536618 357959 536621
rect 399845 536618 399954 536621
rect 357893 536616 360210 536618
rect 357893 536560 357898 536616
rect 357954 536560 360210 536616
rect 357893 536558 360210 536560
rect 399764 536616 399954 536618
rect 399764 536560 399850 536616
rect 399906 536560 399954 536616
rect 399764 536558 399954 536560
rect 357893 536555 357959 536558
rect 322473 536210 322539 536213
rect 319854 536208 322539 536210
rect 319854 536152 322478 536208
rect 322534 536152 322539 536208
rect 319854 536150 322539 536152
rect 322473 536147 322539 536150
rect 360150 536112 360210 536558
rect 399845 536555 399954 536558
rect 399894 536346 399954 536555
rect 400765 536346 400831 536349
rect 399894 536344 400831 536346
rect 399894 536288 400770 536344
rect 400826 536288 400831 536344
rect 399894 536286 400831 536288
rect 400765 536283 400831 536286
rect 401593 536210 401659 536213
rect 399894 536208 401659 536210
rect 399894 536152 401598 536208
rect 401654 536152 401659 536208
rect 399894 536150 401659 536152
rect 399894 536112 399954 536150
rect 401593 536147 401659 536150
rect 399334 535604 399340 535668
rect 399404 535666 399410 535668
rect 399753 535666 399819 535669
rect 399404 535664 399819 535666
rect 399404 535608 399758 535664
rect 399814 535608 399819 535664
rect 399404 535606 399819 535608
rect 399404 535604 399410 535606
rect 399753 535603 399819 535606
rect 400397 535462 400463 535465
rect 399924 535460 400463 535462
rect 254669 535394 254735 535397
rect 322197 535394 322263 535397
rect 251804 535392 254735 535394
rect 251804 535336 254674 535392
rect 254730 535336 254735 535392
rect 251804 535334 254735 535336
rect 254669 535331 254735 535334
rect 319854 535392 322263 535394
rect 319854 535336 322202 535392
rect 322258 535336 322263 535392
rect 319854 535334 322263 535336
rect 319854 535296 319914 535334
rect 322197 535331 322263 535334
rect 357433 535394 357499 535397
rect 360150 535394 360210 535432
rect 399924 535404 400402 535460
rect 400458 535404 400463 535460
rect 399924 535402 400463 535404
rect 400397 535399 400463 535402
rect 357433 535392 360210 535394
rect 357433 535336 357438 535392
rect 357494 535336 360210 535392
rect 357433 535334 360210 535336
rect 357433 535331 357499 535334
rect 357433 534986 357499 534989
rect 357433 534984 360210 534986
rect 357433 534928 357438 534984
rect 357494 534928 360210 534984
rect 357433 534926 360210 534928
rect 357433 534923 357499 534926
rect 360150 534752 360210 534926
rect 401869 534714 401935 534717
rect 399894 534712 401935 534714
rect 399894 534656 401874 534712
rect 401930 534656 401935 534712
rect 399894 534654 401935 534656
rect 319854 534442 319914 534616
rect 357525 534578 357591 534581
rect 357525 534576 360210 534578
rect 357525 534520 357530 534576
rect 357586 534520 360210 534576
rect 357525 534518 360210 534520
rect 357525 534515 357591 534518
rect 322473 534442 322539 534445
rect 319854 534440 322539 534442
rect 319854 534384 322478 534440
rect 322534 534384 322539 534440
rect 319854 534382 322539 534384
rect 322473 534379 322539 534382
rect 360150 534072 360210 534518
rect 399894 534072 399954 534654
rect 401869 534651 401935 534654
rect 322381 534034 322447 534037
rect 319854 534032 322447 534034
rect 319854 533976 322386 534032
rect 322442 533976 322447 534032
rect 319854 533974 322447 533976
rect 319854 533936 319914 533974
rect 322381 533971 322447 533974
rect 401869 533762 401935 533765
rect 399894 533760 401935 533762
rect 399894 533704 401874 533760
rect 401930 533704 401935 533760
rect 399894 533702 401935 533704
rect 399894 533392 399954 533702
rect 401869 533699 401935 533702
rect 322841 533354 322907 533357
rect 319854 533352 322907 533354
rect 319854 533296 322846 533352
rect 322902 533296 322907 533352
rect 319854 533294 322907 533296
rect 319854 533256 319914 533294
rect 322841 533291 322907 533294
rect 357709 533354 357775 533357
rect 360150 533354 360210 533392
rect 357709 533352 360210 533354
rect 357709 533296 357714 533352
rect 357770 533296 360210 533352
rect 357709 533294 360210 533296
rect 357709 533291 357775 533294
rect 399334 533156 399340 533220
rect 399404 533218 399410 533220
rect 399753 533218 399819 533221
rect 401777 533218 401843 533221
rect 399404 533216 399819 533218
rect 399404 533160 399758 533216
rect 399814 533160 399819 533216
rect 399404 533158 399819 533160
rect 399404 533156 399410 533158
rect 399753 533155 399819 533158
rect 399894 533216 401843 533218
rect 399894 533160 401782 533216
rect 401838 533160 401843 533216
rect 399894 533158 401843 533160
rect 358905 532810 358971 532813
rect 358905 532808 360210 532810
rect 358905 532752 358910 532808
rect 358966 532752 360210 532808
rect 358905 532750 360210 532752
rect 358905 532747 358971 532750
rect 360150 532712 360210 532750
rect 399894 532712 399954 533158
rect 401777 533155 401843 533158
rect 481582 532612 481588 532676
rect 481652 532674 481658 532676
rect 481817 532674 481883 532677
rect 481652 532672 481883 532674
rect 481652 532616 481822 532672
rect 481878 532616 481883 532672
rect 481652 532614 481883 532616
rect 481652 532612 481658 532614
rect 481817 532611 481883 532614
rect 484669 532674 484735 532677
rect 484894 532674 484900 532676
rect 484669 532672 484900 532674
rect 484669 532616 484674 532672
rect 484730 532616 484900 532672
rect 484669 532614 484900 532616
rect 484669 532611 484735 532614
rect 484894 532612 484900 532614
rect 484964 532612 484970 532676
rect 488993 532674 489059 532677
rect 489126 532674 489132 532676
rect 488993 532672 489132 532674
rect 488993 532616 488998 532672
rect 489054 532616 489132 532672
rect 488993 532614 489132 532616
rect 488993 532611 489059 532614
rect 489126 532612 489132 532614
rect 489196 532612 489202 532676
rect 501873 532674 501939 532677
rect 502006 532674 502012 532676
rect 501873 532672 502012 532674
rect 501873 532616 501878 532672
rect 501934 532616 502012 532672
rect 501873 532614 502012 532616
rect 501873 532611 501939 532614
rect 502006 532612 502012 532614
rect 502076 532612 502082 532676
rect 50981 532402 51047 532405
rect 319854 532402 319914 532576
rect 402421 532538 402487 532541
rect 399894 532536 402487 532538
rect 399894 532480 402426 532536
rect 402482 532480 402487 532536
rect 399894 532478 402487 532480
rect 322197 532402 322263 532405
rect 50981 532400 52164 532402
rect 50981 532344 50986 532400
rect 51042 532344 52164 532400
rect 50981 532342 52164 532344
rect 319854 532400 322263 532402
rect 319854 532344 322202 532400
rect 322258 532344 322263 532400
rect 319854 532342 322263 532344
rect 50981 532339 51047 532342
rect 322197 532339 322263 532342
rect 357433 532402 357499 532405
rect 357433 532400 360210 532402
rect 357433 532344 357438 532400
rect 357494 532344 360210 532400
rect 357433 532342 360210 532344
rect 357433 532339 357499 532342
rect 321645 532266 321711 532269
rect 319854 532264 321711 532266
rect 319854 532208 321650 532264
rect 321706 532208 321711 532264
rect 319854 532206 321711 532208
rect 319854 531896 319914 532206
rect 321645 532203 321711 532206
rect 360150 532032 360210 532342
rect 399894 532032 399954 532478
rect 402421 532475 402487 532478
rect 499430 532476 499436 532540
rect 499500 532538 499506 532540
rect 500953 532538 501019 532541
rect 499500 532536 501019 532538
rect 499500 532480 500958 532536
rect 501014 532480 501019 532536
rect 499500 532478 501019 532480
rect 499500 532476 499506 532478
rect 500953 532475 501019 532478
rect 357525 531858 357591 531861
rect 401961 531858 402027 531861
rect 357525 531856 360210 531858
rect 357525 531800 357530 531856
rect 357586 531800 360210 531856
rect 357525 531798 360210 531800
rect 357525 531795 357591 531798
rect 360150 531352 360210 531798
rect 399894 531856 402027 531858
rect 399894 531800 401966 531856
rect 402022 531800 402027 531856
rect 399894 531798 402027 531800
rect 399894 531352 399954 531798
rect 401961 531795 402027 531798
rect 319854 531178 319914 531216
rect 322473 531178 322539 531181
rect 319854 531176 322539 531178
rect 319854 531120 322478 531176
rect 322534 531120 322539 531176
rect 319854 531118 322539 531120
rect 322473 531115 322539 531118
rect 330477 530634 330543 530637
rect 353477 530634 353543 530637
rect 358486 530634 358492 530636
rect 330477 530632 358492 530634
rect 330477 530576 330482 530632
rect 330538 530576 353482 530632
rect 353538 530576 358492 530632
rect 330477 530574 358492 530576
rect 330477 530571 330543 530574
rect 353477 530571 353543 530574
rect 358486 530572 358492 530574
rect 358556 530634 358562 530636
rect 358556 530574 360210 530634
rect 358556 530572 358562 530574
rect 319854 530226 319914 530536
rect 322381 530226 322447 530229
rect 319854 530224 322447 530226
rect 319854 530168 322386 530224
rect 322442 530168 322447 530224
rect 319854 530166 322447 530168
rect 322381 530163 322447 530166
rect 360150 529992 360210 530574
rect 399894 530362 399954 530672
rect 402881 530362 402947 530365
rect 399894 530360 402947 530362
rect 399894 530304 402886 530360
rect 402942 530304 402947 530360
rect 399894 530302 402947 530304
rect 402881 530299 402947 530302
rect 401961 530226 402027 530229
rect 399894 530224 402027 530226
rect 399894 530168 401966 530224
rect 402022 530168 402027 530224
rect 399894 530166 402027 530168
rect 399894 529992 399954 530166
rect 401961 530163 402027 530166
rect 482921 529954 482987 529957
rect 484158 529954 484164 529956
rect 482921 529952 484164 529954
rect 482921 529896 482926 529952
rect 482982 529896 484164 529952
rect 482921 529894 484164 529896
rect 482921 529891 482987 529894
rect 484158 529892 484164 529894
rect 484228 529892 484234 529956
rect 319854 529818 319914 529856
rect 322473 529818 322539 529821
rect 319854 529816 322539 529818
rect 319854 529760 322478 529816
rect 322534 529760 322539 529816
rect 319854 529758 322539 529760
rect 322473 529755 322539 529758
rect 477493 529682 477559 529685
rect 477493 529680 480178 529682
rect 477493 529624 477498 529680
rect 477554 529624 480178 529680
rect 477493 529622 480178 529624
rect 477493 529619 477559 529622
rect 254209 529546 254275 529549
rect 251804 529544 254275 529546
rect 251804 529488 254214 529544
rect 254270 529488 254275 529544
rect 251804 529486 254275 529488
rect 254209 529483 254275 529486
rect 357433 529546 357499 529549
rect 357433 529544 360210 529546
rect 357433 529488 357438 529544
rect 357494 529488 360210 529544
rect 357433 529486 360210 529488
rect 357433 529483 357499 529486
rect 360150 529312 360210 529486
rect 480118 529312 480178 529622
rect 489545 529546 489611 529549
rect 502425 529548 502491 529549
rect 489678 529546 489684 529548
rect 489545 529544 489684 529546
rect 489545 529488 489550 529544
rect 489606 529488 489684 529544
rect 489545 529486 489684 529488
rect 489545 529483 489611 529486
rect 489678 529484 489684 529486
rect 489748 529484 489754 529548
rect 502374 529546 502380 529548
rect 502334 529486 502380 529546
rect 502444 529544 502491 529548
rect 502486 529488 502491 529544
rect 502374 529484 502380 529486
rect 502444 529484 502491 529488
rect 503662 529484 503668 529548
rect 503732 529546 503738 529548
rect 504173 529546 504239 529549
rect 503732 529544 504239 529546
rect 503732 529488 504178 529544
rect 504234 529488 504239 529544
rect 503732 529486 504239 529488
rect 503732 529484 503738 529486
rect 502425 529483 502491 529484
rect 504173 529483 504239 529486
rect 319854 528866 319914 529176
rect 399894 529002 399954 529312
rect 402881 529002 402947 529005
rect 399894 529000 402947 529002
rect 399894 528944 402886 529000
rect 402942 528944 402947 529000
rect 399894 528942 402947 528944
rect 509926 529002 509986 529312
rect 511165 529002 511231 529005
rect 509926 529000 511231 529002
rect 509926 528944 511170 529000
rect 511226 528944 511231 529000
rect 509926 528942 511231 528944
rect 402881 528939 402947 528942
rect 511165 528939 511231 528942
rect 322749 528866 322815 528869
rect 403157 528866 403223 528869
rect 319854 528864 322815 528866
rect 319854 528808 322754 528864
rect 322810 528808 322815 528864
rect 319854 528806 322815 528808
rect 322749 528803 322815 528806
rect 399894 528864 403223 528866
rect 399894 528808 403162 528864
rect 403218 528808 403223 528864
rect 399894 528806 403223 528808
rect 399894 528632 399954 528806
rect 403157 528803 403223 528806
rect 358169 528594 358235 528597
rect 360150 528594 360210 528632
rect 358169 528592 360210 528594
rect 358169 528536 358174 528592
rect 358230 528536 360210 528592
rect 358169 528534 360210 528536
rect 477493 528594 477559 528597
rect 480118 528594 480178 528632
rect 477493 528592 480178 528594
rect 477493 528536 477498 528592
rect 477554 528536 480178 528592
rect 477493 528534 480178 528536
rect 509926 528594 509986 528632
rect 513281 528594 513347 528597
rect 509926 528592 513347 528594
rect 509926 528536 513286 528592
rect 513342 528536 513347 528592
rect 509926 528534 513347 528536
rect 358169 528531 358235 528534
rect 477493 528531 477559 528534
rect 513281 528531 513347 528534
rect 319854 528458 319914 528496
rect 322289 528458 322355 528461
rect 402881 528458 402947 528461
rect 319854 528456 322355 528458
rect 319854 528400 322294 528456
rect 322350 528400 322355 528456
rect 319854 528398 322355 528400
rect 322289 528395 322355 528398
rect 399894 528456 402947 528458
rect 399894 528400 402886 528456
rect 402942 528400 402947 528456
rect 399894 528398 402947 528400
rect 359365 528322 359431 528325
rect 359365 528320 360210 528322
rect 359365 528264 359370 528320
rect 359426 528264 360210 528320
rect 359365 528262 360210 528264
rect 359365 528259 359431 528262
rect 322473 528186 322539 528189
rect 319854 528184 322539 528186
rect 319854 528128 322478 528184
rect 322534 528128 322539 528184
rect 319854 528126 322539 528128
rect -960 527764 480 528004
rect 319854 527816 319914 528126
rect 322473 528123 322539 528126
rect 360150 527952 360210 528262
rect 399894 527952 399954 528398
rect 402881 528395 402947 528398
rect 358537 527778 358603 527781
rect 401961 527778 402027 527781
rect 358537 527776 360210 527778
rect 358537 527720 358542 527776
rect 358598 527720 360210 527776
rect 358537 527718 360210 527720
rect 358537 527715 358603 527718
rect 360150 527272 360210 527718
rect 399894 527776 402027 527778
rect 399894 527720 401966 527776
rect 402022 527720 402027 527776
rect 399894 527718 402027 527720
rect 399894 527272 399954 527718
rect 401961 527715 402027 527718
rect 479149 527506 479215 527509
rect 480118 527506 480178 527952
rect 509374 527508 509434 527952
rect 479149 527504 480178 527506
rect 479149 527448 479154 527504
rect 479210 527448 480178 527504
rect 479149 527446 480178 527448
rect 479149 527443 479215 527446
rect 509366 527444 509372 527508
rect 509436 527444 509442 527508
rect 477493 527234 477559 527237
rect 480118 527234 480178 527272
rect 477493 527232 480178 527234
rect 477493 527176 477498 527232
rect 477554 527176 480178 527232
rect 477493 527174 480178 527176
rect 509926 527234 509986 527272
rect 512545 527234 512611 527237
rect 509926 527232 512611 527234
rect 509926 527176 512550 527232
rect 512606 527176 512611 527232
rect 509926 527174 512611 527176
rect 477493 527171 477559 527174
rect 512545 527171 512611 527174
rect 319854 527098 319914 527136
rect 321553 527098 321619 527101
rect 400673 527098 400739 527101
rect 401777 527098 401843 527101
rect 319854 527096 321619 527098
rect 319854 527040 321558 527096
rect 321614 527040 321619 527096
rect 319854 527038 321619 527040
rect 321553 527035 321619 527038
rect 399894 527096 401843 527098
rect 399894 527040 400678 527096
rect 400734 527040 401782 527096
rect 401838 527040 401843 527096
rect 399894 527038 401843 527040
rect 358537 526962 358603 526965
rect 360510 526962 360516 526964
rect 358537 526960 360516 526962
rect 358537 526904 358542 526960
rect 358598 526904 360516 526960
rect 358537 526902 360516 526904
rect 358537 526899 358603 526902
rect 360510 526900 360516 526902
rect 360580 526900 360586 526964
rect 322473 526826 322539 526829
rect 319854 526824 322539 526826
rect 319854 526768 322478 526824
rect 322534 526768 322539 526824
rect 319854 526766 322539 526768
rect 50889 526554 50955 526557
rect 50889 526552 52164 526554
rect 50889 526496 50894 526552
rect 50950 526496 52164 526552
rect 50889 526494 52164 526496
rect 50889 526491 50955 526494
rect 319854 526456 319914 526766
rect 322473 526763 322539 526766
rect 357433 526826 357499 526829
rect 357433 526824 360210 526826
rect 357433 526768 357438 526824
rect 357494 526768 360210 526824
rect 357433 526766 360210 526768
rect 357433 526763 357499 526766
rect 360150 526592 360210 526766
rect 399894 526592 399954 527038
rect 400673 527035 400739 527038
rect 401777 527035 401843 527038
rect 357893 526418 357959 526421
rect 402237 526418 402303 526421
rect 357893 526416 360210 526418
rect 357893 526360 357898 526416
rect 357954 526360 360210 526416
rect 357893 526358 360210 526360
rect 357893 526355 357959 526358
rect 360150 525912 360210 526358
rect 399894 526416 402303 526418
rect 399894 526360 402242 526416
rect 402298 526360 402303 526416
rect 399894 526358 402303 526360
rect 399894 525912 399954 526358
rect 402237 526355 402303 526358
rect 479057 526146 479123 526149
rect 480118 526146 480178 526592
rect 509926 526554 509986 526592
rect 510613 526554 510679 526557
rect 511073 526554 511139 526557
rect 509926 526552 511139 526554
rect 509926 526496 510618 526552
rect 510674 526496 511078 526552
rect 511134 526496 511139 526552
rect 509926 526494 511139 526496
rect 510613 526491 510679 526494
rect 511073 526491 511139 526494
rect 512269 526418 512335 526421
rect 479057 526144 480178 526146
rect 479057 526088 479062 526144
rect 479118 526088 480178 526144
rect 479057 526086 480178 526088
rect 509926 526416 512335 526418
rect 509926 526360 512274 526416
rect 512330 526360 512335 526416
rect 509926 526358 512335 526360
rect 479057 526083 479123 526086
rect 509926 525912 509986 526358
rect 512269 526355 512335 526358
rect 477493 525874 477559 525877
rect 480118 525874 480178 525912
rect 477493 525872 480178 525874
rect 477493 525816 477498 525872
rect 477554 525816 480178 525872
rect 477493 525814 480178 525816
rect 477493 525811 477559 525814
rect 319854 525738 319914 525776
rect 322473 525738 322539 525741
rect 319854 525736 322539 525738
rect 319854 525680 322478 525736
rect 322534 525680 322539 525736
rect 319854 525678 322539 525680
rect 322473 525675 322539 525678
rect 477953 525602 478019 525605
rect 477953 525600 480178 525602
rect 477953 525544 477958 525600
rect 478014 525544 480178 525600
rect 477953 525542 480178 525544
rect 477953 525539 478019 525542
rect 400305 525262 400371 525265
rect 399924 525260 400371 525262
rect 358077 525194 358143 525197
rect 360150 525194 360210 525232
rect 399924 525204 400310 525260
rect 400366 525204 400371 525260
rect 480118 525232 480178 525542
rect 399924 525202 400371 525204
rect 400305 525199 400371 525202
rect 358077 525192 360210 525194
rect 358077 525136 358082 525192
rect 358138 525136 360210 525192
rect 358077 525134 360210 525136
rect 358077 525131 358143 525134
rect 319854 524650 319914 525096
rect 358629 525058 358695 525061
rect 402237 525058 402303 525061
rect 358629 525056 360210 525058
rect 358629 525000 358634 525056
rect 358690 525000 360210 525056
rect 358629 524998 360210 525000
rect 358629 524995 358695 524998
rect 322565 524650 322631 524653
rect 319854 524648 322631 524650
rect 319854 524592 322570 524648
rect 322626 524592 322631 524648
rect 319854 524590 322631 524592
rect 322565 524587 322631 524590
rect 360150 524552 360210 524998
rect 399894 525056 402303 525058
rect 399894 525000 402242 525056
rect 402298 525000 402303 525056
rect 399894 524998 402303 525000
rect 399894 524552 399954 524998
rect 402237 524995 402303 524998
rect 478689 525058 478755 525061
rect 478689 525056 480178 525058
rect 478689 525000 478694 525056
rect 478750 525000 480178 525056
rect 478689 524998 480178 525000
rect 478689 524995 478755 524998
rect 480118 524552 480178 524998
rect 509926 524922 509986 525232
rect 512637 524922 512703 524925
rect 509926 524920 512703 524922
rect 509926 524864 512642 524920
rect 512698 524864 512703 524920
rect 509926 524862 512703 524864
rect 512637 524859 512703 524862
rect 322289 524514 322355 524517
rect 319854 524512 322355 524514
rect 319854 524456 322294 524512
rect 322350 524456 322355 524512
rect 319854 524454 322355 524456
rect 509926 524514 509986 524552
rect 512361 524514 512427 524517
rect 509926 524512 512427 524514
rect 509926 524456 512366 524512
rect 512422 524456 512427 524512
rect 509926 524454 512427 524456
rect 319854 524416 319914 524454
rect 322289 524451 322355 524454
rect 512361 524451 512427 524454
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 402881 524106 402947 524109
rect 399894 524104 402947 524106
rect 399894 524048 402886 524104
rect 402942 524048 402947 524104
rect 399894 524046 402947 524048
rect 399894 523872 399954 524046
rect 402881 524043 402947 524046
rect 358629 523834 358695 523837
rect 360150 523834 360210 523872
rect 358629 523832 360210 523834
rect 358629 523776 358634 523832
rect 358690 523776 360210 523832
rect 358629 523774 360210 523776
rect 358629 523771 358695 523774
rect 254025 523698 254091 523701
rect 251804 523696 254091 523698
rect 251804 523640 254030 523696
rect 254086 523640 254091 523696
rect 251804 523638 254091 523640
rect 254025 523635 254091 523638
rect 319854 523426 319914 523736
rect 357433 523698 357499 523701
rect 399569 523698 399635 523701
rect 357433 523696 360210 523698
rect 357433 523640 357438 523696
rect 357494 523640 360210 523696
rect 357433 523638 360210 523640
rect 357433 523635 357499 523638
rect 322473 523426 322539 523429
rect 319854 523424 322539 523426
rect 319854 523368 322478 523424
rect 322534 523368 322539 523424
rect 319854 523366 322539 523368
rect 322473 523363 322539 523366
rect 360150 523192 360210 523638
rect 399526 523696 399635 523698
rect 399526 523640 399574 523696
rect 399630 523640 399635 523696
rect 399526 523635 399635 523640
rect 399526 523192 399586 523635
rect 477493 523426 477559 523429
rect 480118 523426 480178 523872
rect 477493 523424 480178 523426
rect 477493 523368 477498 523424
rect 477554 523368 480178 523424
rect 477493 523366 480178 523368
rect 509926 523426 509986 523872
rect 512545 523426 512611 523429
rect 509926 523424 512611 523426
rect 509926 523368 512550 523424
rect 512606 523368 512611 523424
rect 509926 523366 512611 523368
rect 477493 523363 477559 523366
rect 512545 523363 512611 523366
rect 322381 523154 322447 523157
rect 319854 523152 322447 523154
rect 319854 523096 322386 523152
rect 322442 523096 322447 523152
rect 319854 523094 322447 523096
rect 319854 523056 319914 523094
rect 322381 523091 322447 523094
rect 477493 523154 477559 523157
rect 480118 523154 480178 523192
rect 477493 523152 480178 523154
rect 477493 523096 477498 523152
rect 477554 523096 480178 523152
rect 477493 523094 480178 523096
rect 477493 523091 477559 523094
rect 509926 523021 509986 523192
rect 400489 523018 400555 523021
rect 399894 523016 400555 523018
rect 399894 522960 400494 523016
rect 400550 522960 400555 523016
rect 399894 522958 400555 522960
rect 399894 522512 399954 522958
rect 400489 522955 400555 522958
rect 509877 523016 509986 523021
rect 509877 522960 509882 523016
rect 509938 522960 509986 523016
rect 509877 522958 509986 522960
rect 509877 522955 509943 522958
rect 319854 522066 319914 522376
rect 322473 522066 322539 522069
rect 319854 522064 322539 522066
rect 319854 522008 322478 522064
rect 322534 522008 322539 522064
rect 319854 522006 322539 522008
rect 322473 522003 322539 522006
rect 358445 522066 358511 522069
rect 360150 522066 360210 522512
rect 358445 522064 360210 522066
rect 358445 522008 358450 522064
rect 358506 522008 360210 522064
rect 358445 522006 360210 522008
rect 478413 522066 478479 522069
rect 480118 522066 480178 522512
rect 478413 522064 480178 522066
rect 478413 522008 478418 522064
rect 478474 522008 480178 522064
rect 478413 522006 480178 522008
rect 509926 522066 509986 522512
rect 512453 522066 512519 522069
rect 509926 522064 512519 522066
rect 509926 522008 512458 522064
rect 512514 522008 512519 522064
rect 509926 522006 512519 522008
rect 358445 522003 358511 522006
rect 478413 522003 478479 522006
rect 512453 522003 512519 522006
rect 322013 521930 322079 521933
rect 319854 521928 322079 521930
rect 319854 521872 322018 521928
rect 322074 521872 322079 521928
rect 319854 521870 322079 521872
rect 319854 521696 319914 521870
rect 322013 521867 322079 521870
rect 357985 521930 358051 521933
rect 357985 521928 360210 521930
rect 357985 521872 357990 521928
rect 358046 521872 360210 521928
rect 357985 521870 360210 521872
rect 357985 521867 358051 521870
rect 360150 521832 360210 521870
rect 399894 521794 399954 521832
rect 402881 521794 402947 521797
rect 399894 521792 402947 521794
rect 399894 521736 402886 521792
rect 402942 521736 402947 521792
rect 399894 521734 402947 521736
rect 402881 521731 402947 521734
rect 477953 521794 478019 521797
rect 480118 521794 480178 521832
rect 477953 521792 480178 521794
rect 477953 521736 477958 521792
rect 478014 521736 480178 521792
rect 477953 521734 480178 521736
rect 509926 521794 509986 521832
rect 512821 521794 512887 521797
rect 509926 521792 512887 521794
rect 509926 521736 512826 521792
rect 512882 521736 512887 521792
rect 509926 521734 512887 521736
rect 477953 521731 478019 521734
rect 512821 521731 512887 521734
rect 49325 521660 49391 521661
rect 49325 521658 49372 521660
rect 49280 521656 49372 521658
rect 49280 521600 49330 521656
rect 49280 521598 49372 521600
rect 49325 521596 49372 521598
rect 49436 521596 49442 521660
rect 359089 521658 359155 521661
rect 359089 521656 360210 521658
rect 359089 521600 359094 521656
rect 359150 521600 360210 521656
rect 359089 521598 360210 521600
rect 49325 521595 49391 521596
rect 359089 521595 359155 521598
rect 360150 521152 360210 521598
rect 399334 521596 399340 521660
rect 399404 521596 399410 521660
rect 399342 521152 399402 521596
rect 49325 520706 49391 520709
rect 319854 520706 319914 521016
rect 359273 520978 359339 520981
rect 401593 520978 401659 520981
rect 359273 520976 360210 520978
rect 359273 520920 359278 520976
rect 359334 520920 360210 520976
rect 359273 520918 360210 520920
rect 359273 520915 359339 520918
rect 322473 520706 322539 520709
rect 49325 520704 52164 520706
rect 49325 520648 49330 520704
rect 49386 520648 52164 520704
rect 49325 520646 52164 520648
rect 319854 520704 322539 520706
rect 319854 520648 322478 520704
rect 322534 520648 322539 520704
rect 319854 520646 322539 520648
rect 49325 520643 49391 520646
rect 322473 520643 322539 520646
rect 322013 520570 322079 520573
rect 319854 520568 322079 520570
rect 319854 520512 322018 520568
rect 322074 520512 322079 520568
rect 319854 520510 322079 520512
rect 319854 520336 319914 520510
rect 322013 520507 322079 520510
rect 360150 520472 360210 520918
rect 399894 520976 401659 520978
rect 399894 520920 401598 520976
rect 401654 520920 401659 520976
rect 399894 520918 401659 520920
rect 399894 520472 399954 520918
rect 401593 520915 401659 520918
rect 477493 520706 477559 520709
rect 480118 520706 480178 521152
rect 477493 520704 480178 520706
rect 477493 520648 477498 520704
rect 477554 520648 480178 520704
rect 477493 520646 480178 520648
rect 509926 520706 509986 521152
rect 512913 520706 512979 520709
rect 509926 520704 512979 520706
rect 509926 520648 512918 520704
rect 512974 520648 512979 520704
rect 509926 520646 512979 520648
rect 477493 520643 477559 520646
rect 512913 520643 512979 520646
rect 478597 520298 478663 520301
rect 480118 520298 480178 520472
rect 478597 520296 480178 520298
rect 478597 520240 478602 520296
rect 478658 520240 480178 520296
rect 478597 520238 480178 520240
rect 509926 520298 509986 520472
rect 510981 520298 511047 520301
rect 509926 520296 511047 520298
rect 509926 520240 510986 520296
rect 511042 520240 511047 520296
rect 509926 520238 511047 520240
rect 478597 520235 478663 520238
rect 510981 520235 511047 520238
rect 401593 520162 401659 520165
rect 399894 520160 401659 520162
rect 399894 520104 401598 520160
rect 401654 520104 401659 520160
rect 399894 520102 401659 520104
rect 399894 519792 399954 520102
rect 401593 520099 401659 520102
rect 358261 519754 358327 519757
rect 360150 519754 360210 519792
rect 358261 519752 360210 519754
rect 358261 519696 358266 519752
rect 358322 519696 360210 519752
rect 358261 519694 360210 519696
rect 358261 519691 358327 519694
rect 319854 519346 319914 519656
rect 357433 519618 357499 519621
rect 357433 519616 360210 519618
rect 357433 519560 357438 519616
rect 357494 519560 360210 519616
rect 357433 519558 360210 519560
rect 357433 519555 357499 519558
rect 321553 519346 321619 519349
rect 319854 519344 321619 519346
rect 319854 519288 321558 519344
rect 321614 519288 321619 519344
rect 319854 519286 321619 519288
rect 321553 519283 321619 519286
rect 322841 519210 322907 519213
rect 319854 519208 322907 519210
rect 319854 519152 322846 519208
rect 322902 519152 322907 519208
rect 319854 519150 322907 519152
rect 319854 518976 319914 519150
rect 322841 519147 322907 519150
rect 360150 519112 360210 519558
rect 478505 519346 478571 519349
rect 480118 519346 480178 519792
rect 478505 519344 480178 519346
rect 478505 519288 478510 519344
rect 478566 519288 480178 519344
rect 478505 519286 480178 519288
rect 509926 519346 509986 519792
rect 510797 519346 510863 519349
rect 509926 519344 510863 519346
rect 509926 519288 510802 519344
rect 510858 519288 510863 519344
rect 509926 519286 510863 519288
rect 478505 519283 478571 519286
rect 510797 519283 510863 519286
rect 478689 519074 478755 519077
rect 480118 519074 480178 519112
rect 478689 519072 480178 519074
rect 478689 519016 478694 519072
rect 478750 519016 480178 519072
rect 478689 519014 480178 519016
rect 509926 519074 509986 519112
rect 513281 519074 513347 519077
rect 509926 519072 513347 519074
rect 509926 519016 513286 519072
rect 513342 519016 513347 519072
rect 509926 519014 513347 519016
rect 478689 519011 478755 519014
rect 513281 519011 513347 519014
rect 325693 518938 325759 518941
rect 326981 518938 327047 518941
rect 349102 518938 349108 518940
rect 325693 518936 349108 518938
rect 325693 518880 325698 518936
rect 325754 518880 326986 518936
rect 327042 518880 349108 518936
rect 325693 518878 349108 518880
rect 325693 518875 325759 518878
rect 326981 518875 327047 518878
rect 349102 518876 349108 518878
rect 349172 518876 349178 518940
rect 357433 518802 357499 518805
rect 357433 518800 360210 518802
rect 357433 518744 357438 518800
rect 357494 518744 360210 518800
rect 357433 518742 360210 518744
rect 357433 518739 357499 518742
rect 360150 518432 360210 518742
rect 399334 518740 399340 518804
rect 399404 518740 399410 518804
rect 399342 518432 399402 518740
rect 319854 517986 319914 518296
rect 402513 518258 402579 518261
rect 399894 518256 402579 518258
rect 399894 518200 402518 518256
rect 402574 518200 402579 518256
rect 399894 518198 402579 518200
rect 322473 517986 322539 517989
rect 319854 517984 322539 517986
rect 319854 517928 322478 517984
rect 322534 517928 322539 517984
rect 319854 517926 322539 517928
rect 322473 517923 322539 517926
rect 254485 517850 254551 517853
rect 321829 517850 321895 517853
rect 251804 517848 254551 517850
rect 251804 517792 254490 517848
rect 254546 517792 254551 517848
rect 251804 517790 254551 517792
rect 254485 517787 254551 517790
rect 319854 517848 321895 517850
rect 319854 517792 321834 517848
rect 321890 517792 321895 517848
rect 319854 517790 321895 517792
rect 319854 517616 319914 517790
rect 321829 517787 321895 517790
rect 399894 517752 399954 518198
rect 402513 518195 402579 518198
rect 477585 517986 477651 517989
rect 480118 517986 480178 518432
rect 477585 517984 480178 517986
rect 477585 517928 477590 517984
rect 477646 517928 480178 517984
rect 477585 517926 480178 517928
rect 509742 517989 509802 518432
rect 512177 518258 512243 518261
rect 509926 518256 512243 518258
rect 509926 518200 512182 518256
rect 512238 518200 512243 518256
rect 509926 518198 512243 518200
rect 509742 517984 509851 517989
rect 509742 517928 509790 517984
rect 509846 517928 509851 517984
rect 509742 517926 509851 517928
rect 477585 517923 477651 517926
rect 509785 517923 509851 517926
rect 509926 517752 509986 518198
rect 512177 518195 512243 518198
rect 357525 517578 357591 517581
rect 360150 517578 360210 517752
rect 477493 517714 477559 517717
rect 480118 517714 480178 517752
rect 477493 517712 480178 517714
rect 477493 517656 477498 517712
rect 477554 517656 480178 517712
rect 477493 517654 480178 517656
rect 477493 517651 477559 517654
rect 357525 517576 360210 517578
rect 357525 517520 357530 517576
rect 357586 517520 360210 517576
rect 357525 517518 360210 517520
rect 357525 517515 357591 517518
rect 321553 517442 321619 517445
rect 319854 517440 321619 517442
rect 319854 517384 321558 517440
rect 321614 517384 321619 517440
rect 319854 517382 321619 517384
rect 319854 516936 319914 517382
rect 321553 517379 321619 517382
rect 357433 517442 357499 517445
rect 402053 517442 402119 517445
rect 357433 517440 360210 517442
rect 357433 517384 357438 517440
rect 357494 517384 360210 517440
rect 357433 517382 360210 517384
rect 357433 517379 357499 517382
rect 360150 517072 360210 517382
rect 399894 517440 402119 517442
rect 399894 517384 402058 517440
rect 402114 517384 402119 517440
rect 399894 517382 402119 517384
rect 399894 517072 399954 517382
rect 402053 517379 402119 517382
rect 478229 517034 478295 517037
rect 480118 517034 480178 517072
rect 478229 517032 480178 517034
rect 478229 516976 478234 517032
rect 478290 516976 480178 517032
rect 478229 516974 480178 516976
rect 478229 516971 478295 516974
rect 478505 516898 478571 516901
rect 478505 516896 480178 516898
rect 478505 516840 478510 516896
rect 478566 516840 480178 516896
rect 478505 516838 480178 516840
rect 478505 516835 478571 516838
rect 480118 516392 480178 516838
rect 509926 516626 509986 517072
rect 513189 516626 513255 516629
rect 509926 516624 513255 516626
rect 509926 516568 513194 516624
rect 513250 516568 513255 516624
rect 509926 516566 513255 516568
rect 513189 516563 513255 516566
rect 322381 516354 322447 516357
rect 319854 516352 322447 516354
rect 319854 516296 322386 516352
rect 322442 516296 322447 516352
rect 319854 516294 322447 516296
rect 319854 516256 319914 516294
rect 322381 516291 322447 516294
rect 357157 516218 357223 516221
rect 358537 516218 358603 516221
rect 360150 516218 360210 516392
rect 357157 516216 360210 516218
rect 357157 516160 357162 516216
rect 357218 516160 358542 516216
rect 358598 516160 360210 516216
rect 357157 516158 360210 516160
rect 399894 516218 399954 516392
rect 509926 516354 509986 516392
rect 513281 516354 513347 516357
rect 509926 516352 513347 516354
rect 509926 516296 513286 516352
rect 513342 516296 513347 516352
rect 509926 516294 513347 516296
rect 513281 516291 513347 516294
rect 402605 516218 402671 516221
rect 399894 516216 402671 516218
rect 399894 516160 402610 516216
rect 402666 516160 402671 516216
rect 399894 516158 402671 516160
rect 357157 516155 357223 516158
rect 358537 516155 358603 516158
rect 402605 516155 402671 516158
rect 401593 516082 401659 516085
rect 399894 516080 401659 516082
rect 399894 516024 401598 516080
rect 401654 516024 401659 516080
rect 399894 516022 401659 516024
rect 399894 515712 399954 516022
rect 401593 516019 401659 516022
rect 319854 515538 319914 515576
rect 322841 515538 322907 515541
rect 319854 515536 322907 515538
rect 319854 515480 322846 515536
rect 322902 515480 322907 515536
rect 319854 515478 322907 515480
rect 322841 515475 322907 515478
rect 321829 515402 321895 515405
rect 319854 515400 321895 515402
rect 319854 515344 321834 515400
rect 321890 515344 321895 515400
rect 319854 515342 321895 515344
rect -960 514858 480 514948
rect 319854 514896 319914 515342
rect 321829 515339 321895 515342
rect 358537 515130 358603 515133
rect 360150 515130 360210 515712
rect 400581 515538 400647 515541
rect 401961 515538 402027 515541
rect 358537 515128 360210 515130
rect 358537 515072 358542 515128
rect 358598 515072 360210 515128
rect 358537 515070 360210 515072
rect 399894 515536 402027 515538
rect 399894 515480 400586 515536
rect 400642 515480 401966 515536
rect 402022 515480 402027 515536
rect 399894 515478 402027 515480
rect 358537 515067 358603 515070
rect 399894 515032 399954 515478
rect 400581 515475 400647 515478
rect 401961 515475 402027 515478
rect 478965 515266 479031 515269
rect 480118 515266 480178 515712
rect 509926 515674 509986 515712
rect 512269 515674 512335 515677
rect 509926 515672 512335 515674
rect 509926 515616 512274 515672
rect 512330 515616 512335 515672
rect 509926 515614 512335 515616
rect 512269 515611 512335 515614
rect 513189 515538 513255 515541
rect 478965 515264 480178 515266
rect 478965 515208 478970 515264
rect 479026 515208 480178 515264
rect 478965 515206 480178 515208
rect 509926 515536 513255 515538
rect 509926 515480 513194 515536
rect 513250 515480 513255 515536
rect 509926 515478 513255 515480
rect 478965 515203 479031 515206
rect 509926 515032 509986 515478
rect 513189 515475 513255 515478
rect 3693 514858 3759 514861
rect -960 514856 3759 514858
rect -960 514800 3698 514856
rect 3754 514800 3759 514856
rect -960 514798 3759 514800
rect -960 514708 480 514798
rect 3693 514795 3759 514798
rect 51073 514858 51139 514861
rect 479241 514858 479307 514861
rect 480118 514858 480178 515032
rect 51073 514856 52164 514858
rect 51073 514800 51078 514856
rect 51134 514800 52164 514856
rect 51073 514798 52164 514800
rect 479241 514856 480178 514858
rect 479241 514800 479246 514856
rect 479302 514800 480178 514856
rect 479241 514798 480178 514800
rect 51073 514795 51139 514798
rect 479241 514795 479307 514798
rect 357433 514722 357499 514725
rect 357433 514720 360210 514722
rect 357433 514664 357438 514720
rect 357494 514664 360210 514720
rect 357433 514662 360210 514664
rect 357433 514659 357499 514662
rect 360150 514352 360210 514662
rect 510981 514450 511047 514453
rect 509926 514448 511047 514450
rect 509926 514392 510986 514448
rect 511042 514392 511047 514448
rect 509926 514390 511047 514392
rect 509926 514352 509986 514390
rect 510981 514387 511047 514390
rect 319854 514178 319914 514216
rect 321645 514178 321711 514181
rect 322105 514178 322171 514181
rect 319854 514176 322171 514178
rect 319854 514120 321650 514176
rect 321706 514120 322110 514176
rect 322166 514120 322171 514176
rect 319854 514118 322171 514120
rect 321645 514115 321711 514118
rect 322105 514115 322171 514118
rect 399894 513906 399954 514352
rect 401593 513906 401659 513909
rect 399894 513904 401659 513906
rect 399894 513848 401598 513904
rect 401654 513848 401659 513904
rect 399894 513846 401659 513848
rect 401593 513843 401659 513846
rect 477585 513906 477651 513909
rect 480118 513906 480178 514352
rect 510705 514314 510771 514317
rect 510110 514312 510771 514314
rect 510110 514256 510710 514312
rect 510766 514256 510771 514312
rect 510110 514254 510771 514256
rect 510110 514178 510170 514254
rect 510705 514251 510771 514254
rect 477585 513904 480178 513906
rect 477585 513848 477590 513904
rect 477646 513848 480178 513904
rect 477585 513846 480178 513848
rect 509926 514118 510170 514178
rect 477585 513843 477651 513846
rect 509926 513672 509986 514118
rect 319854 513498 319914 513536
rect 322473 513498 322539 513501
rect 360150 513498 360210 513672
rect 319854 513496 322539 513498
rect 319854 513440 322478 513496
rect 322534 513440 322539 513496
rect 319854 513438 322539 513440
rect 322473 513435 322539 513438
rect 358310 513438 360210 513498
rect 399894 513498 399954 513672
rect 402053 513498 402119 513501
rect 399894 513496 402119 513498
rect 399894 513440 402058 513496
rect 402114 513440 402119 513496
rect 399894 513438 402119 513440
rect 358310 513229 358370 513438
rect 402053 513435 402119 513438
rect 477493 513498 477559 513501
rect 480118 513498 480178 513672
rect 477493 513496 480178 513498
rect 477493 513440 477498 513496
rect 477554 513440 480178 513496
rect 477493 513438 480178 513440
rect 477493 513435 477559 513438
rect 358997 513362 359063 513365
rect 358997 513360 360210 513362
rect 358997 513304 359002 513360
rect 359058 513304 360210 513360
rect 358997 513302 360210 513304
rect 358997 513299 359063 513302
rect 358261 513224 358370 513229
rect 358261 513168 358266 513224
rect 358322 513168 358370 513224
rect 358261 513166 358370 513168
rect 358261 513163 358327 513166
rect 360150 512992 360210 513302
rect 402513 513226 402579 513229
rect 399894 513224 402579 513226
rect 399894 513168 402518 513224
rect 402574 513168 402579 513224
rect 399894 513166 402579 513168
rect 399894 512992 399954 513166
rect 402513 513163 402579 513166
rect 510061 513022 510127 513025
rect 509956 513020 510127 513022
rect 478781 512954 478847 512957
rect 480118 512954 480178 512992
rect 509956 512964 510066 513020
rect 510122 512964 510127 513020
rect 509956 512962 510127 512964
rect 510061 512959 510127 512962
rect 478781 512952 480178 512954
rect 478781 512896 478786 512952
rect 478842 512896 480178 512952
rect 478781 512894 480178 512896
rect 478781 512891 478847 512894
rect 319854 512682 319914 512856
rect 357433 512818 357499 512821
rect 402421 512818 402487 512821
rect 357433 512816 360210 512818
rect 357433 512760 357438 512816
rect 357494 512760 360210 512816
rect 357433 512758 360210 512760
rect 357433 512755 357499 512758
rect 321737 512682 321803 512685
rect 322105 512682 322171 512685
rect 319854 512680 322171 512682
rect 319854 512624 321742 512680
rect 321798 512624 322110 512680
rect 322166 512624 322171 512680
rect 319854 512622 322171 512624
rect 321737 512619 321803 512622
rect 322105 512619 322171 512622
rect 360150 512312 360210 512758
rect 399894 512816 402487 512818
rect 399894 512760 402426 512816
rect 402482 512760 402487 512816
rect 399894 512758 402487 512760
rect 399894 512312 399954 512758
rect 402421 512755 402487 512758
rect 477585 512818 477651 512821
rect 512126 512818 512132 512820
rect 477585 512816 480178 512818
rect 477585 512760 477590 512816
rect 477646 512760 480178 512816
rect 477585 512758 480178 512760
rect 477585 512755 477651 512758
rect 480118 512312 480178 512758
rect 509926 512758 512132 512818
rect 509926 512312 509986 512758
rect 512126 512756 512132 512758
rect 512196 512756 512202 512820
rect 320357 512206 320423 512209
rect 319884 512204 320466 512206
rect 319884 512148 320362 512204
rect 320418 512148 320466 512204
rect 319884 512146 320466 512148
rect 320357 512143 320466 512146
rect 320406 512138 320466 512143
rect 320909 512138 320975 512141
rect 320406 512136 320975 512138
rect 320406 512080 320914 512136
rect 320970 512080 320975 512136
rect 320406 512078 320975 512080
rect 320909 512075 320975 512078
rect 254393 512002 254459 512005
rect 402329 512002 402395 512005
rect 251804 512000 254459 512002
rect 251804 511944 254398 512000
rect 254454 511944 254459 512000
rect 251804 511942 254459 511944
rect 254393 511939 254459 511942
rect 399894 512000 402395 512002
rect 399894 511944 402334 512000
rect 402390 511944 402395 512000
rect 399894 511942 402395 511944
rect 399894 511632 399954 511942
rect 402329 511939 402395 511942
rect 357617 511594 357683 511597
rect 360150 511594 360210 511632
rect 357617 511592 360210 511594
rect 357617 511536 357622 511592
rect 357678 511536 360210 511592
rect 357617 511534 360210 511536
rect 357617 511531 357683 511534
rect 319854 511322 319914 511496
rect 357433 511458 357499 511461
rect 357433 511456 360210 511458
rect 357433 511400 357438 511456
rect 357494 511400 360210 511456
rect 357433 511398 360210 511400
rect 357433 511395 357499 511398
rect 321553 511322 321619 511325
rect 319854 511320 321619 511322
rect 319854 511264 321558 511320
rect 321614 511264 321619 511320
rect 319854 511262 321619 511264
rect 321553 511259 321619 511262
rect 360150 510952 360210 511398
rect 477585 511186 477651 511189
rect 480118 511186 480178 511632
rect 477585 511184 480178 511186
rect 477585 511128 477590 511184
rect 477646 511128 480178 511184
rect 477585 511126 480178 511128
rect 509926 511189 509986 511632
rect 580349 511322 580415 511325
rect 583520 511322 584960 511412
rect 580349 511320 584960 511322
rect 580349 511264 580354 511320
rect 580410 511264 584960 511320
rect 580349 511262 584960 511264
rect 580349 511259 580415 511262
rect 509926 511184 510035 511189
rect 509926 511128 509974 511184
rect 510030 511128 510035 511184
rect 583520 511172 584960 511262
rect 509926 511126 510035 511128
rect 477585 511123 477651 511126
rect 509969 511123 510035 511126
rect 320357 510846 320423 510849
rect 319884 510844 320423 510846
rect 319884 510788 320362 510844
rect 320418 510788 320423 510844
rect 319884 510786 320423 510788
rect 320357 510783 320423 510786
rect 399894 510778 399954 510952
rect 402881 510778 402947 510781
rect 399894 510776 402947 510778
rect 399894 510720 402886 510776
rect 402942 510720 402947 510776
rect 399894 510718 402947 510720
rect 402881 510715 402947 510718
rect 477861 510642 477927 510645
rect 480118 510642 480178 510952
rect 509926 510778 509986 510952
rect 513281 510778 513347 510781
rect 509926 510776 513347 510778
rect 509926 510720 513286 510776
rect 513342 510720 513347 510776
rect 509926 510718 513347 510720
rect 513281 510715 513347 510718
rect 477861 510640 480178 510642
rect 477861 510584 477866 510640
rect 477922 510584 480178 510640
rect 477861 510582 480178 510584
rect 477861 510579 477927 510582
rect 401869 510506 401935 510509
rect 399894 510504 401935 510506
rect 399894 510448 401874 510504
rect 401930 510448 401935 510504
rect 399894 510446 401935 510448
rect 357433 510370 357499 510373
rect 357433 510368 360210 510370
rect 357433 510312 357438 510368
rect 357494 510312 360210 510368
rect 357433 510310 360210 510312
rect 357433 510307 357499 510310
rect 360150 510272 360210 510310
rect 399894 510272 399954 510446
rect 401869 510443 401935 510446
rect 477493 510506 477559 510509
rect 477493 510504 480178 510506
rect 477493 510448 477498 510504
rect 477554 510448 480178 510504
rect 477493 510446 480178 510448
rect 477493 510443 477559 510446
rect 480118 510272 480178 510446
rect 510429 510302 510495 510305
rect 509956 510300 510495 510302
rect 509956 510244 510434 510300
rect 510490 510244 510495 510300
rect 509956 510242 510495 510244
rect 510429 510239 510495 510242
rect 320081 510166 320147 510169
rect 319884 510164 320147 510166
rect 319884 510136 320086 510164
rect 319854 510108 320086 510136
rect 320142 510108 320147 510164
rect 319854 510106 320147 510108
rect 319345 509962 319411 509965
rect 319854 509962 319914 510106
rect 320081 510103 320147 510106
rect 357801 510098 357867 510101
rect 357801 510096 360210 510098
rect 357801 510040 357806 510096
rect 357862 510040 360210 510096
rect 357801 510038 360210 510040
rect 357801 510035 357867 510038
rect 319345 509960 319914 509962
rect 319345 509904 319350 509960
rect 319406 509904 319914 509960
rect 319345 509902 319914 509904
rect 319345 509899 319411 509902
rect 360150 509592 360210 510038
rect 320449 509554 320515 509557
rect 319854 509552 320515 509554
rect 319854 509496 320454 509552
rect 320510 509496 320515 509552
rect 319854 509494 320515 509496
rect 399894 509554 399954 509592
rect 402881 509554 402947 509557
rect 399894 509552 402947 509554
rect 399894 509496 402886 509552
rect 402942 509496 402947 509552
rect 399894 509494 402947 509496
rect 319854 509456 319914 509494
rect 320449 509491 320515 509494
rect 402881 509491 402947 509494
rect 404905 509420 404971 509421
rect 404854 509418 404860 509420
rect 404814 509358 404860 509418
rect 404924 509416 404971 509420
rect 404966 509360 404971 509416
rect 404854 509356 404860 509358
rect 404924 509356 404971 509360
rect 404905 509355 404971 509356
rect 477493 509418 477559 509421
rect 480118 509418 480178 509592
rect 477493 509416 480178 509418
rect 477493 509360 477498 509416
rect 477554 509360 480178 509416
rect 477493 509358 480178 509360
rect 509926 509418 509986 509592
rect 513281 509418 513347 509421
rect 509926 509416 513347 509418
rect 509926 509360 513286 509416
rect 513342 509360 513347 509416
rect 509926 509358 513347 509360
rect 477493 509355 477559 509358
rect 513281 509355 513347 509358
rect 50797 509010 50863 509013
rect 357433 509010 357499 509013
rect 50797 509008 52164 509010
rect 50797 508952 50802 509008
rect 50858 508952 52164 509008
rect 50797 508950 52164 508952
rect 357433 509008 360210 509010
rect 357433 508952 357438 509008
rect 357494 508952 360210 509008
rect 357433 508950 360210 508952
rect 50797 508947 50863 508950
rect 357433 508947 357499 508950
rect 360150 508912 360210 508950
rect 319302 508333 319362 508776
rect 357525 508738 357591 508741
rect 357525 508736 360210 508738
rect 357525 508680 357530 508736
rect 357586 508680 360210 508736
rect 357525 508678 360210 508680
rect 357525 508675 357591 508678
rect 319302 508328 319411 508333
rect 319302 508272 319350 508328
rect 319406 508272 319411 508328
rect 319302 508270 319411 508272
rect 319345 508267 319411 508270
rect 360150 508232 360210 508678
rect 399894 508466 399954 508912
rect 401869 508466 401935 508469
rect 480118 508466 480178 508912
rect 399894 508464 401935 508466
rect 399894 508408 401874 508464
rect 401930 508408 401935 508464
rect 399894 508406 401935 508408
rect 401869 508403 401935 508406
rect 479750 508406 480178 508466
rect 401726 508330 401732 508332
rect 399894 508270 401732 508330
rect 399894 508232 399954 508270
rect 401726 508268 401732 508270
rect 401796 508268 401802 508332
rect 478781 508330 478847 508333
rect 479750 508330 479810 508406
rect 478781 508328 479810 508330
rect 478781 508272 478786 508328
rect 478842 508272 479810 508328
rect 478781 508270 479810 508272
rect 478781 508267 478847 508270
rect 320173 508126 320239 508129
rect 319884 508124 320466 508126
rect 319884 508068 320178 508124
rect 320234 508068 320466 508124
rect 319884 508066 320466 508068
rect 320173 508063 320239 508066
rect 320406 508058 320466 508066
rect 320541 508058 320607 508061
rect 320406 508056 320607 508058
rect 320406 508000 320546 508056
rect 320602 508000 320607 508056
rect 320406 507998 320607 508000
rect 320541 507995 320607 507998
rect 478505 507922 478571 507925
rect 480118 507922 480178 508232
rect 478505 507920 480178 507922
rect 478505 507864 478510 507920
rect 478566 507864 480178 507920
rect 478505 507862 480178 507864
rect 509926 507922 509986 508232
rect 511257 507922 511323 507925
rect 509926 507920 511323 507922
rect 509926 507864 511262 507920
rect 511318 507864 511323 507920
rect 509926 507862 511323 507864
rect 478505 507859 478571 507862
rect 511257 507859 511323 507862
rect 357801 507786 357867 507789
rect 357801 507784 360210 507786
rect 357801 507728 357806 507784
rect 357862 507728 360210 507784
rect 357801 507726 360210 507728
rect 357801 507723 357867 507726
rect 360150 507552 360210 507726
rect 399334 507724 399340 507788
rect 399404 507724 399410 507788
rect 399342 507552 399402 507724
rect 320357 507446 320423 507449
rect 319884 507444 320423 507446
rect 319884 507388 320362 507444
rect 320418 507388 320423 507444
rect 319884 507386 320423 507388
rect 320357 507383 320423 507386
rect 357433 507378 357499 507381
rect 399477 507378 399543 507381
rect 357433 507376 360210 507378
rect 357433 507320 357438 507376
rect 357494 507320 360210 507376
rect 357433 507318 360210 507320
rect 357433 507315 357499 507318
rect 360150 506872 360210 507318
rect 399477 507376 399586 507378
rect 399477 507320 399482 507376
rect 399538 507320 399586 507376
rect 399477 507315 399586 507320
rect 399526 506872 399586 507315
rect 478137 507106 478203 507109
rect 480118 507106 480178 507552
rect 478137 507104 480178 507106
rect 478137 507048 478142 507104
rect 478198 507048 480178 507104
rect 478137 507046 480178 507048
rect 509926 507106 509986 507552
rect 510705 507106 510771 507109
rect 509926 507104 510771 507106
rect 509926 507048 510710 507104
rect 510766 507048 510771 507104
rect 509926 507046 510771 507048
rect 478137 507043 478203 507046
rect 510705 507043 510771 507046
rect 320081 506766 320147 506769
rect 319884 506764 320147 506766
rect 319884 506708 320086 506764
rect 320142 506708 320147 506764
rect 319884 506706 320147 506708
rect 320081 506703 320147 506706
rect 479425 506562 479491 506565
rect 480118 506562 480178 506872
rect 479425 506560 480178 506562
rect 479425 506504 479430 506560
rect 479486 506504 480178 506560
rect 479425 506502 480178 506504
rect 509926 506562 509986 506872
rect 512913 506562 512979 506565
rect 509926 506560 512979 506562
rect 509926 506504 512918 506560
rect 512974 506504 512979 506560
rect 509926 506502 512979 506504
rect 479425 506499 479491 506502
rect 512913 506499 512979 506502
rect 402237 506426 402303 506429
rect 399894 506424 402303 506426
rect 399894 506368 402242 506424
rect 402298 506368 402303 506424
rect 399894 506366 402303 506368
rect 357433 506290 357499 506293
rect 357433 506288 360210 506290
rect 357433 506232 357438 506288
rect 357494 506232 360210 506288
rect 357433 506230 360210 506232
rect 357433 506227 357499 506230
rect 360150 506192 360210 506230
rect 399894 506192 399954 506366
rect 402237 506363 402303 506366
rect 254301 506154 254367 506157
rect 251804 506152 254367 506154
rect 251804 506096 254306 506152
rect 254362 506096 254367 506152
rect 251804 506094 254367 506096
rect 254301 506091 254367 506094
rect 319302 505613 319362 506056
rect 402145 506018 402211 506021
rect 399894 506016 402211 506018
rect 399894 505960 402150 506016
rect 402206 505960 402211 506016
rect 399894 505958 402211 505960
rect 357525 505882 357591 505885
rect 357525 505880 360210 505882
rect 357525 505824 357530 505880
rect 357586 505824 360210 505880
rect 357525 505822 360210 505824
rect 357525 505819 357591 505822
rect 319302 505608 319411 505613
rect 319302 505552 319350 505608
rect 319406 505552 319411 505608
rect 319302 505550 319411 505552
rect 319345 505547 319411 505550
rect 360150 505512 360210 505822
rect 399894 505512 399954 505958
rect 402145 505955 402211 505958
rect 477493 505746 477559 505749
rect 480118 505746 480178 506192
rect 477493 505744 480178 505746
rect 477493 505688 477498 505744
rect 477554 505688 480178 505744
rect 477493 505686 480178 505688
rect 509926 505746 509986 506192
rect 510981 505746 511047 505749
rect 509926 505744 511047 505746
rect 509926 505688 510986 505744
rect 511042 505688 511047 505744
rect 509926 505686 511047 505688
rect 477493 505683 477559 505686
rect 510981 505683 511047 505686
rect 510245 505542 510311 505545
rect 509956 505540 510311 505542
rect 320173 505406 320239 505409
rect 319884 505404 320239 505406
rect 319884 505348 320178 505404
rect 320234 505348 320239 505404
rect 319884 505346 320239 505348
rect 320173 505343 320239 505346
rect 477493 505338 477559 505341
rect 480118 505338 480178 505512
rect 509956 505484 510250 505540
rect 510306 505484 510311 505540
rect 509956 505482 510311 505484
rect 510245 505479 510311 505482
rect 477493 505336 480178 505338
rect 477493 505280 477498 505336
rect 477554 505280 480178 505336
rect 477493 505278 480178 505280
rect 477493 505275 477559 505278
rect 358854 505004 358860 505068
rect 358924 505066 358930 505068
rect 358924 505006 360210 505066
rect 358924 505004 358930 505006
rect 360150 504832 360210 505006
rect 400438 504862 400444 504864
rect 399924 504802 400444 504862
rect 400438 504800 400444 504802
rect 400508 504800 400514 504864
rect 320081 504726 320147 504729
rect 319884 504724 320147 504726
rect 319884 504696 320086 504724
rect 319854 504668 320086 504696
rect 320142 504668 320147 504724
rect 319854 504666 320147 504668
rect 319345 504250 319411 504253
rect 319854 504250 319914 504666
rect 320081 504663 320147 504666
rect 357433 504658 357499 504661
rect 357433 504656 360210 504658
rect 357433 504600 357438 504656
rect 357494 504600 360210 504656
rect 357433 504598 360210 504600
rect 357433 504595 357499 504598
rect 319345 504248 319914 504250
rect 319345 504192 319350 504248
rect 319406 504192 319914 504248
rect 319345 504190 319914 504192
rect 319345 504187 319411 504190
rect 360150 504152 360210 504598
rect 477585 504386 477651 504389
rect 480118 504386 480178 504832
rect 477585 504384 480178 504386
rect 477585 504328 477590 504384
rect 477646 504328 480178 504384
rect 477585 504326 480178 504328
rect 509926 504386 509986 504832
rect 511349 504386 511415 504389
rect 509926 504384 511415 504386
rect 509926 504328 511354 504384
rect 511410 504328 511415 504384
rect 509926 504326 511415 504328
rect 477585 504323 477651 504326
rect 511349 504323 511415 504326
rect 400213 504182 400279 504185
rect 399924 504180 400279 504182
rect 399924 504124 400218 504180
rect 400274 504124 400279 504180
rect 399924 504122 400279 504124
rect 400213 504119 400279 504122
rect 322381 504114 322447 504117
rect 319854 504112 322447 504114
rect 319854 504056 322386 504112
rect 322442 504056 322447 504112
rect 319854 504054 322447 504056
rect 319854 504016 319914 504054
rect 322381 504051 322447 504054
rect 477493 503978 477559 503981
rect 480118 503978 480178 504152
rect 477493 503976 480178 503978
rect 477493 503920 477498 503976
rect 477554 503920 480178 503976
rect 477493 503918 480178 503920
rect 509926 503978 509986 504152
rect 513281 503978 513347 503981
rect 509926 503976 513347 503978
rect 509926 503920 513286 503976
rect 513342 503920 513347 503976
rect 509926 503918 513347 503920
rect 477493 503915 477559 503918
rect 513281 503915 513347 503918
rect 358721 503706 358787 503709
rect 511993 503706 512059 503709
rect 358721 503704 360210 503706
rect 358721 503648 358726 503704
rect 358782 503648 360210 503704
rect 358721 503646 360210 503648
rect 358721 503643 358787 503646
rect 360150 503472 360210 503646
rect 509926 503704 512059 503706
rect 509926 503648 511998 503704
rect 512054 503648 512059 503704
rect 509926 503646 512059 503648
rect 509926 503472 509986 503646
rect 511993 503643 512059 503646
rect 322381 503434 322447 503437
rect 319854 503432 322447 503434
rect 319854 503376 322386 503432
rect 322442 503376 322447 503432
rect 319854 503374 322447 503376
rect 319854 503336 319914 503374
rect 322381 503371 322447 503374
rect 357433 503298 357499 503301
rect 401685 503298 401751 503301
rect 357433 503296 360210 503298
rect 357433 503240 357438 503296
rect 357494 503240 360210 503296
rect 357433 503238 360210 503240
rect 357433 503235 357499 503238
rect 49233 503162 49299 503165
rect 49550 503162 49556 503164
rect 49233 503160 49556 503162
rect 49233 503104 49238 503160
rect 49294 503104 49556 503160
rect 49233 503102 49556 503104
rect 49233 503099 49299 503102
rect 49550 503100 49556 503102
rect 49620 503162 49626 503164
rect 49620 503102 52164 503162
rect 49620 503100 49626 503102
rect 360150 502792 360210 503238
rect 399894 503296 401751 503298
rect 399894 503240 401690 503296
rect 401746 503240 401751 503296
rect 399894 503238 401751 503240
rect 399894 502792 399954 503238
rect 401685 503235 401751 503238
rect 479333 503026 479399 503029
rect 480118 503026 480178 503472
rect 479333 503024 480178 503026
rect 479333 502968 479338 503024
rect 479394 502968 480178 503024
rect 479333 502966 480178 502968
rect 479333 502963 479399 502966
rect 319854 502482 319914 502656
rect 477493 502618 477559 502621
rect 480118 502618 480178 502792
rect 477493 502616 480178 502618
rect 477493 502560 477498 502616
rect 477554 502560 480178 502616
rect 477493 502558 480178 502560
rect 509926 502618 509986 502792
rect 513281 502618 513347 502621
rect 509926 502616 513347 502618
rect 509926 502560 513286 502616
rect 513342 502560 513347 502616
rect 509926 502558 513347 502560
rect 477493 502555 477559 502558
rect 513281 502555 513347 502558
rect 322381 502482 322447 502485
rect 319854 502480 322447 502482
rect 319854 502424 322386 502480
rect 322442 502424 322447 502480
rect 319854 502422 322447 502424
rect 322381 502419 322447 502422
rect 358670 502284 358676 502348
rect 358740 502346 358746 502348
rect 358740 502286 360210 502346
rect 358740 502284 358746 502286
rect 360150 502112 360210 502286
rect 510337 502142 510403 502145
rect 509956 502140 510403 502142
rect 357433 501938 357499 501941
rect 357433 501936 360210 501938
rect -960 501802 480 501892
rect 357433 501880 357438 501936
rect 357494 501880 360210 501936
rect 357433 501878 360210 501880
rect 357433 501875 357499 501878
rect 3601 501802 3667 501805
rect -960 501800 3667 501802
rect -960 501744 3606 501800
rect 3662 501744 3667 501800
rect -960 501742 3667 501744
rect -960 501652 480 501742
rect 3601 501739 3667 501742
rect 360150 501432 360210 501878
rect 399526 501669 399586 502112
rect 399477 501664 399586 501669
rect 399477 501608 399482 501664
rect 399538 501608 399586 501664
rect 399477 501606 399586 501608
rect 477493 501666 477559 501669
rect 480118 501666 480178 502112
rect 509956 502084 510342 502140
rect 510398 502084 510403 502140
rect 509956 502082 510403 502084
rect 510337 502079 510403 502082
rect 477493 501664 480178 501666
rect 477493 501608 477498 501664
rect 477554 501608 480178 501664
rect 477493 501606 480178 501608
rect 399477 501603 399543 501606
rect 477493 501603 477559 501606
rect 400254 501462 400260 501464
rect 399924 501402 400260 501462
rect 400254 501400 400260 501402
rect 400324 501400 400330 501464
rect 359406 501196 359412 501260
rect 359476 501258 359482 501260
rect 359476 501198 360210 501258
rect 359476 501196 359482 501198
rect 360150 500752 360210 501198
rect 478781 500986 478847 500989
rect 480118 500986 480178 501432
rect 478781 500984 480178 500986
rect 478781 500928 478786 500984
rect 478842 500928 480178 500984
rect 478781 500926 480178 500928
rect 509926 500986 509986 501432
rect 511993 500986 512059 500989
rect 509926 500984 512059 500986
rect 509926 500928 511998 500984
rect 512054 500928 512059 500984
rect 509926 500926 512059 500928
rect 478781 500923 478847 500926
rect 511993 500923 512059 500926
rect 512085 500850 512151 500853
rect 509926 500848 512151 500850
rect 509926 500792 512090 500848
rect 512146 500792 512151 500848
rect 509926 500790 512151 500792
rect 509926 500752 509986 500790
rect 512085 500787 512151 500790
rect 254209 500306 254275 500309
rect 251804 500304 254275 500306
rect 251804 500248 254214 500304
rect 254270 500248 254275 500304
rect 251804 500246 254275 500248
rect 399894 500306 399954 500752
rect 401869 500306 401935 500309
rect 399894 500304 401935 500306
rect 399894 500248 401874 500304
rect 401930 500248 401935 500304
rect 399894 500246 401935 500248
rect 254209 500243 254275 500246
rect 401869 500243 401935 500246
rect 477493 500170 477559 500173
rect 480118 500170 480178 500752
rect 477493 500168 480178 500170
rect 477493 500112 477498 500168
rect 477554 500112 480178 500168
rect 477493 500110 480178 500112
rect 477493 500107 477559 500110
rect 360653 499898 360719 499901
rect 361430 499898 361436 499900
rect 360653 499896 361436 499898
rect 360653 499840 360658 499896
rect 360714 499840 361436 499896
rect 360653 499838 361436 499840
rect 360653 499835 360719 499838
rect 361430 499836 361436 499838
rect 361500 499836 361506 499900
rect 361614 499836 361620 499900
rect 361684 499898 361690 499900
rect 362585 499898 362651 499901
rect 361684 499896 362651 499898
rect 361684 499840 362590 499896
rect 362646 499840 362651 499896
rect 361684 499838 362651 499840
rect 361684 499836 361690 499838
rect 362585 499835 362651 499838
rect 364742 499836 364748 499900
rect 364812 499898 364818 499900
rect 365161 499898 365227 499901
rect 364812 499896 365227 499898
rect 364812 499840 365166 499896
rect 365222 499840 365227 499896
rect 364812 499838 365227 499840
rect 364812 499836 364818 499838
rect 365161 499835 365227 499838
rect 368238 499836 368244 499900
rect 368308 499898 368314 499900
rect 368381 499898 368447 499901
rect 368308 499896 368447 499898
rect 368308 499840 368386 499896
rect 368442 499840 368447 499896
rect 368308 499838 368447 499840
rect 368308 499836 368314 499838
rect 368381 499835 368447 499838
rect 368606 499836 368612 499900
rect 368676 499898 368682 499900
rect 369669 499898 369735 499901
rect 368676 499896 369735 499898
rect 368676 499840 369674 499896
rect 369730 499840 369735 499896
rect 368676 499838 369735 499840
rect 368676 499836 368682 499838
rect 369669 499835 369735 499838
rect 370078 499836 370084 499900
rect 370148 499898 370154 499900
rect 370313 499898 370379 499901
rect 370148 499896 370379 499898
rect 370148 499840 370318 499896
rect 370374 499840 370379 499896
rect 370148 499838 370379 499840
rect 370148 499836 370154 499838
rect 370313 499835 370379 499838
rect 373758 499836 373764 499900
rect 373828 499898 373834 499900
rect 374821 499898 374887 499901
rect 373828 499896 374887 499898
rect 373828 499840 374826 499896
rect 374882 499840 374887 499896
rect 373828 499838 374887 499840
rect 373828 499836 373834 499838
rect 374821 499835 374887 499838
rect 376109 499898 376175 499901
rect 376334 499898 376340 499900
rect 376109 499896 376340 499898
rect 376109 499840 376114 499896
rect 376170 499840 376340 499896
rect 376109 499838 376340 499840
rect 376109 499835 376175 499838
rect 376334 499836 376340 499838
rect 376404 499836 376410 499900
rect 376753 499898 376819 499901
rect 380617 499900 380683 499901
rect 376886 499898 376892 499900
rect 376753 499896 376892 499898
rect 376753 499840 376758 499896
rect 376814 499840 376892 499896
rect 376753 499838 376892 499840
rect 376753 499835 376819 499838
rect 376886 499836 376892 499838
rect 376956 499836 376962 499900
rect 380566 499836 380572 499900
rect 380636 499898 380683 499900
rect 380636 499896 380728 499898
rect 380678 499840 380728 499896
rect 380636 499838 380728 499840
rect 380636 499836 380683 499838
rect 380934 499836 380940 499900
rect 381004 499898 381010 499900
rect 381261 499898 381327 499901
rect 381004 499896 381327 499898
rect 381004 499840 381266 499896
rect 381322 499840 381327 499896
rect 381004 499838 381327 499840
rect 381004 499836 381010 499838
rect 380617 499835 380683 499836
rect 381261 499835 381327 499838
rect 382549 499898 382615 499901
rect 382774 499898 382780 499900
rect 382549 499896 382780 499898
rect 382549 499840 382554 499896
rect 382610 499840 382780 499896
rect 382549 499838 382780 499840
rect 382549 499835 382615 499838
rect 382774 499836 382780 499838
rect 382844 499836 382850 499900
rect 385125 499898 385191 499901
rect 385534 499898 385540 499900
rect 385125 499896 385540 499898
rect 385125 499840 385130 499896
rect 385186 499840 385540 499896
rect 385125 499838 385540 499840
rect 385125 499835 385191 499838
rect 385534 499836 385540 499838
rect 385604 499836 385610 499900
rect 389582 499836 389588 499900
rect 389652 499898 389658 499900
rect 390277 499898 390343 499901
rect 389652 499896 390343 499898
rect 389652 499840 390282 499896
rect 390338 499840 390343 499896
rect 389652 499838 390343 499840
rect 389652 499836 389658 499838
rect 390277 499835 390343 499838
rect 391974 499836 391980 499900
rect 392044 499898 392050 499900
rect 392853 499898 392919 499901
rect 392044 499896 392919 499898
rect 392044 499840 392858 499896
rect 392914 499840 392919 499896
rect 392044 499838 392919 499840
rect 392044 499836 392050 499838
rect 392853 499835 392919 499838
rect 396574 499836 396580 499900
rect 396644 499898 396650 499900
rect 398649 499898 398715 499901
rect 396644 499896 398715 499898
rect 396644 499840 398654 499896
rect 398710 499840 398715 499896
rect 396644 499838 398715 499840
rect 396644 499836 396650 499838
rect 398649 499835 398715 499838
rect 391565 499762 391631 499765
rect 392526 499762 392532 499764
rect 391565 499760 392532 499762
rect 391565 499704 391570 499760
rect 391626 499704 392532 499760
rect 391565 499702 392532 499704
rect 391565 499699 391631 499702
rect 392526 499700 392532 499702
rect 392596 499700 392602 499764
rect 398598 499700 398604 499764
rect 398668 499762 398674 499764
rect 399342 499762 399402 500072
rect 495382 499836 495388 499900
rect 495452 499898 495458 499900
rect 496123 499898 496189 499901
rect 495452 499896 496189 499898
rect 495452 499840 496128 499896
rect 496184 499840 496189 499896
rect 495452 499838 496189 499840
rect 509926 499898 509986 500072
rect 512729 499898 512795 499901
rect 509926 499896 512795 499898
rect 509926 499840 512734 499896
rect 512790 499840 512795 499896
rect 509926 499838 512795 499840
rect 495452 499836 495458 499838
rect 496123 499835 496189 499838
rect 512729 499835 512795 499838
rect 398668 499702 399402 499762
rect 398668 499700 398674 499702
rect 391054 499564 391060 499628
rect 391124 499626 391130 499628
rect 393497 499626 393563 499629
rect 391124 499624 393563 499626
rect 391124 499568 393502 499624
rect 393558 499568 393563 499624
rect 391124 499566 393563 499568
rect 391124 499564 391130 499566
rect 393497 499563 393563 499566
rect 357157 499490 357223 499493
rect 365805 499490 365871 499493
rect 366214 499490 366220 499492
rect 357157 499488 366220 499490
rect 357157 499432 357162 499488
rect 357218 499432 365810 499488
rect 365866 499432 366220 499488
rect 357157 499430 366220 499432
rect 357157 499427 357223 499430
rect 365805 499427 365871 499430
rect 366214 499428 366220 499430
rect 366284 499428 366290 499492
rect 367737 499490 367803 499493
rect 373206 499490 373212 499492
rect 367737 499488 373212 499490
rect 367737 499432 367742 499488
rect 367798 499432 373212 499488
rect 367737 499430 373212 499432
rect 367737 499427 367803 499430
rect 373206 499428 373212 499430
rect 373276 499428 373282 499492
rect 376150 499428 376156 499492
rect 376220 499490 376226 499492
rect 377397 499490 377463 499493
rect 376220 499488 377463 499490
rect 376220 499432 377402 499488
rect 377458 499432 377463 499488
rect 376220 499430 377463 499432
rect 376220 499428 376226 499430
rect 377397 499427 377463 499430
rect 350073 499354 350139 499357
rect 401777 499354 401843 499357
rect 350073 499352 401843 499354
rect 350073 499296 350078 499352
rect 350134 499296 401782 499352
rect 401838 499296 401843 499352
rect 350073 499294 401843 499296
rect 350073 499291 350139 499294
rect 401777 499291 401843 499294
rect 301998 499156 302004 499220
rect 302068 499218 302074 499220
rect 361941 499218 362007 499221
rect 302068 499216 362007 499218
rect 302068 499160 361946 499216
rect 362002 499160 362007 499216
rect 302068 499158 362007 499160
rect 302068 499156 302074 499158
rect 361941 499155 362007 499158
rect 355225 498946 355291 498949
rect 369894 498946 369900 498948
rect 355225 498944 369900 498946
rect 355225 498888 355230 498944
rect 355286 498888 369900 498944
rect 355225 498886 369900 498888
rect 355225 498883 355291 498886
rect 369894 498884 369900 498886
rect 369964 498946 369970 498948
rect 371601 498946 371667 498949
rect 369964 498944 371667 498946
rect 369964 498888 371606 498944
rect 371662 498888 371667 498944
rect 369964 498886 371667 498888
rect 369964 498884 369970 498886
rect 371601 498883 371667 498886
rect 296069 498810 296135 498813
rect 502374 498810 502380 498812
rect 296069 498808 502380 498810
rect 296069 498752 296074 498808
rect 296130 498752 502380 498808
rect 296069 498750 502380 498752
rect 296069 498747 296135 498750
rect 502374 498748 502380 498750
rect 502444 498748 502450 498812
rect 349654 498204 349660 498268
rect 349724 498266 349730 498268
rect 350073 498266 350139 498269
rect 349724 498264 350139 498266
rect 349724 498208 350078 498264
rect 350134 498208 350139 498264
rect 349724 498206 350139 498208
rect 349724 498204 349730 498206
rect 350073 498203 350139 498206
rect 360009 498130 360075 498133
rect 362534 498130 362540 498132
rect 360009 498128 362540 498130
rect 360009 498072 360014 498128
rect 360070 498072 362540 498128
rect 360009 498070 362540 498072
rect 360009 498067 360075 498070
rect 362534 498068 362540 498070
rect 362604 498068 362610 498132
rect 384062 498068 384068 498132
rect 384132 498130 384138 498132
rect 387057 498130 387123 498133
rect 384132 498128 387123 498130
rect 384132 498072 387062 498128
rect 387118 498072 387123 498128
rect 384132 498070 387123 498072
rect 384132 498068 384138 498070
rect 387057 498067 387123 498070
rect 388294 498068 388300 498132
rect 388364 498130 388370 498132
rect 395429 498130 395495 498133
rect 388364 498128 395495 498130
rect 388364 498072 395434 498128
rect 395490 498072 395495 498128
rect 388364 498070 395495 498072
rect 388364 498068 388370 498070
rect 395429 498067 395495 498070
rect 351453 497994 351519 497997
rect 369025 497994 369091 497997
rect 371734 497994 371740 497996
rect 351453 497992 371740 497994
rect 351453 497936 351458 497992
rect 351514 497936 369030 497992
rect 369086 497936 371740 497992
rect 351453 497934 371740 497936
rect 351453 497931 351519 497934
rect 369025 497931 369091 497934
rect 371734 497932 371740 497934
rect 371804 497932 371810 497996
rect 379278 497932 379284 497996
rect 379348 497994 379354 497996
rect 387701 497994 387767 497997
rect 379348 497992 387767 497994
rect 379348 497936 387706 497992
rect 387762 497936 387767 497992
rect 379348 497934 387767 497936
rect 379348 497932 379354 497934
rect 387701 497931 387767 497934
rect 355501 497858 355567 497861
rect 362902 497858 362908 497860
rect 355501 497856 362908 497858
rect 355501 497800 355506 497856
rect 355562 497800 362908 497856
rect 355501 497798 362908 497800
rect 355501 497795 355567 497798
rect 362902 497796 362908 497798
rect 362972 497858 362978 497860
rect 363873 497858 363939 497861
rect 362972 497856 363939 497858
rect 362972 497800 363878 497856
rect 363934 497800 363939 497856
rect 362972 497798 363939 497800
rect 362972 497796 362978 497798
rect 363873 497795 363939 497798
rect 364057 497858 364123 497861
rect 385125 497858 385191 497861
rect 364057 497856 385191 497858
rect 364057 497800 364062 497856
rect 364118 497800 385130 497856
rect 385186 497800 385191 497856
rect 583520 497844 584960 498084
rect 364057 497798 385191 497800
rect 364057 497795 364123 497798
rect 385125 497795 385191 497798
rect 362953 497722 363019 497725
rect 385769 497722 385835 497725
rect 387006 497722 387012 497724
rect 362953 497720 387012 497722
rect 362953 497664 362958 497720
rect 363014 497664 385774 497720
rect 385830 497664 387012 497720
rect 362953 497662 387012 497664
rect 362953 497659 363019 497662
rect 385769 497659 385835 497662
rect 387006 497660 387012 497662
rect 387076 497660 387082 497724
rect 349889 497586 349955 497589
rect 382549 497586 382615 497589
rect 349889 497584 382615 497586
rect 349889 497528 349894 497584
rect 349950 497528 382554 497584
rect 382610 497528 382615 497584
rect 349889 497526 382615 497528
rect 349889 497523 349955 497526
rect 382549 497523 382615 497526
rect 355869 497450 355935 497453
rect 364057 497450 364123 497453
rect 376109 497450 376175 497453
rect 355869 497448 364123 497450
rect 355869 497392 355874 497448
rect 355930 497392 364062 497448
rect 364118 497392 364123 497448
rect 355869 497390 364123 497392
rect 355869 497387 355935 497390
rect 364057 497387 364123 497390
rect 364290 497448 376175 497450
rect 364290 497392 376114 497448
rect 376170 497392 376175 497448
rect 364290 497390 376175 497392
rect 49601 497314 49667 497317
rect 356881 497314 356947 497317
rect 364290 497314 364350 497390
rect 376109 497387 376175 497390
rect 49601 497312 52164 497314
rect 49601 497256 49606 497312
rect 49662 497256 52164 497312
rect 49601 497254 52164 497256
rect 356881 497312 364350 497314
rect 356881 497256 356886 497312
rect 356942 497256 364350 497312
rect 356881 497254 364350 497256
rect 49601 497251 49667 497254
rect 356881 497251 356947 497254
rect 373390 497252 373396 497316
rect 373460 497314 373466 497316
rect 386413 497314 386479 497317
rect 373460 497312 386479 497314
rect 373460 497256 386418 497312
rect 386474 497256 386479 497312
rect 373460 497254 386479 497256
rect 373460 497252 373466 497254
rect 386413 497251 386479 497254
rect 360837 497178 360903 497181
rect 391565 497178 391631 497181
rect 360837 497176 391631 497178
rect 360837 497120 360842 497176
rect 360898 497120 391570 497176
rect 391626 497120 391631 497176
rect 360837 497118 391631 497120
rect 360837 497115 360903 497118
rect 391565 497115 391631 497118
rect 48865 496906 48931 496909
rect 49601 496906 49667 496909
rect 48865 496904 49667 496906
rect 48865 496848 48870 496904
rect 48926 496848 49606 496904
rect 49662 496848 49667 496904
rect 48865 496846 49667 496848
rect 48865 496843 48931 496846
rect 49601 496843 49667 496846
rect 254577 494458 254643 494461
rect 251804 494456 254643 494458
rect 251804 494400 254582 494456
rect 254638 494400 254643 494456
rect 251804 494398 254643 494400
rect 254577 494395 254643 494398
rect 49509 491466 49575 491469
rect 49509 491464 52164 491466
rect 49509 491408 49514 491464
rect 49570 491408 52164 491464
rect 49509 491406 52164 491408
rect 49509 491403 49575 491406
rect -960 488596 480 488836
rect 254669 488610 254735 488613
rect 251804 488608 254735 488610
rect 251804 488552 254674 488608
rect 254730 488552 254735 488608
rect 251804 488550 254735 488552
rect 254669 488547 254735 488550
rect 51257 485618 51323 485621
rect 51257 485616 52164 485618
rect 51257 485560 51262 485616
rect 51318 485560 52164 485616
rect 51257 485558 52164 485560
rect 51257 485555 51323 485558
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 49550 484332 49556 484396
rect 49620 484394 49626 484396
rect 51257 484394 51323 484397
rect 49620 484392 51323 484394
rect 49620 484336 51262 484392
rect 51318 484336 51323 484392
rect 49620 484334 51323 484336
rect 49620 484332 49626 484334
rect 51257 484331 51323 484334
rect 254393 482762 254459 482765
rect 251804 482760 254459 482762
rect 251804 482704 254398 482760
rect 254454 482704 254459 482760
rect 251804 482702 254459 482704
rect 254393 482699 254459 482702
rect 51206 479708 51212 479772
rect 51276 479770 51282 479772
rect 51276 479710 52164 479770
rect 51276 479708 51282 479710
rect 49366 477532 49372 477596
rect 49436 477594 49442 477596
rect 51206 477594 51212 477596
rect 49436 477534 51212 477594
rect 49436 477532 49442 477534
rect 51206 477532 51212 477534
rect 51276 477532 51282 477596
rect 254209 476914 254275 476917
rect 251804 476912 254275 476914
rect 251804 476856 254214 476912
rect 254270 476856 254275 476912
rect 251804 476854 254275 476856
rect 254209 476851 254275 476854
rect -960 475540 480 475780
rect 48957 473922 49023 473925
rect 48957 473920 52164 473922
rect 48957 473864 48962 473920
rect 49018 473864 52164 473920
rect 48957 473862 52164 473864
rect 48957 473859 49023 473862
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect 254485 471066 254551 471069
rect 251804 471064 254551 471066
rect 251804 471008 254490 471064
rect 254546 471008 254551 471064
rect 251804 471006 254551 471008
rect 254485 471003 254551 471006
rect 48773 468074 48839 468077
rect 48773 468072 52164 468074
rect 48773 468016 48778 468072
rect 48834 468016 52164 468072
rect 48773 468014 52164 468016
rect 48773 468011 48839 468014
rect 254669 465218 254735 465221
rect 251804 465216 254735 465218
rect 251804 465160 254674 465216
rect 254730 465160 254735 465216
rect 251804 465158 254735 465160
rect 254669 465155 254735 465158
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 50797 462226 50863 462229
rect 50797 462224 52164 462226
rect 50797 462168 50802 462224
rect 50858 462168 52164 462224
rect 50797 462166 52164 462168
rect 50797 462163 50863 462166
rect 254301 459370 254367 459373
rect 251804 459368 254367 459370
rect 251804 459312 254306 459368
rect 254362 459312 254367 459368
rect 251804 459310 254367 459312
rect 254301 459307 254367 459310
rect 580441 458146 580507 458149
rect 583520 458146 584960 458236
rect 580441 458144 584960 458146
rect 580441 458088 580446 458144
rect 580502 458088 584960 458144
rect 580441 458086 584960 458088
rect 580441 458083 580507 458086
rect 583520 457996 584960 458086
rect 49785 456378 49851 456381
rect 50705 456378 50771 456381
rect 49785 456376 52164 456378
rect 49785 456320 49790 456376
rect 49846 456320 50710 456376
rect 50766 456320 52164 456376
rect 49785 456318 52164 456320
rect 49785 456315 49851 456318
rect 50705 456315 50771 456318
rect 254669 453522 254735 453525
rect 251804 453520 254735 453522
rect 251804 453464 254674 453520
rect 254730 453464 254735 453520
rect 251804 453462 254735 453464
rect 254669 453459 254735 453462
rect 51257 450530 51323 450533
rect 51257 450528 52164 450530
rect 51257 450472 51262 450528
rect 51318 450472 52164 450528
rect 51257 450470 52164 450472
rect 51257 450467 51323 450470
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 254669 447674 254735 447677
rect 251804 447672 254735 447674
rect 251804 447616 254674 447672
rect 254730 447616 254735 447672
rect 251804 447614 254735 447616
rect 254669 447611 254735 447614
rect 48313 444682 48379 444685
rect 48313 444680 52164 444682
rect 48313 444624 48318 444680
rect 48374 444624 52164 444680
rect 583520 444668 584960 444908
rect 48313 444622 52164 444624
rect 48313 444619 48379 444622
rect 254393 441826 254459 441829
rect 251804 441824 254459 441826
rect 251804 441768 254398 441824
rect 254454 441768 254459 441824
rect 251804 441766 254459 441768
rect 254393 441763 254459 441766
rect 48313 438834 48379 438837
rect 48313 438832 52164 438834
rect 48313 438776 48318 438832
rect 48374 438776 52164 438832
rect 48313 438774 52164 438776
rect 48313 438771 48379 438774
rect -960 436508 480 436748
rect 254669 435978 254735 435981
rect 251804 435976 254735 435978
rect 251804 435920 254674 435976
rect 254730 435920 254735 435976
rect 251804 435918 254735 435920
rect 254669 435915 254735 435918
rect 49141 432986 49207 432989
rect 49141 432984 52164 432986
rect 49141 432928 49146 432984
rect 49202 432928 52164 432984
rect 49141 432926 52164 432928
rect 49141 432923 49207 432926
rect 579613 431626 579679 431629
rect 583520 431626 584960 431716
rect 579613 431624 584960 431626
rect 579613 431568 579618 431624
rect 579674 431568 584960 431624
rect 579613 431566 584960 431568
rect 579613 431563 579679 431566
rect 583520 431476 584960 431566
rect 254209 430130 254275 430133
rect 251804 430128 254275 430130
rect 251804 430072 254214 430128
rect 254270 430072 254275 430128
rect 251804 430070 254275 430072
rect 254209 430067 254275 430070
rect 49417 427138 49483 427141
rect 49417 427136 52164 427138
rect 49417 427080 49422 427136
rect 49478 427080 52164 427136
rect 49417 427078 52164 427080
rect 49417 427075 49483 427078
rect 254669 424282 254735 424285
rect 251804 424280 254735 424282
rect 251804 424224 254674 424280
rect 254730 424224 254735 424280
rect 251804 424222 254735 424224
rect 254669 424219 254735 424222
rect -960 423452 480 423692
rect 47945 421290 48011 421293
rect 47945 421288 52164 421290
rect 47945 421232 47950 421288
rect 48006 421232 52164 421288
rect 47945 421230 52164 421232
rect 47945 421227 48011 421230
rect 254393 418434 254459 418437
rect 251804 418432 254459 418434
rect 251804 418376 254398 418432
rect 254454 418376 254459 418432
rect 251804 418374 254459 418376
rect 254393 418371 254459 418374
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 48037 415442 48103 415445
rect 48037 415440 52164 415442
rect 48037 415384 48042 415440
rect 48098 415384 52164 415440
rect 48037 415382 52164 415384
rect 48037 415379 48103 415382
rect 254669 412586 254735 412589
rect 251804 412584 254735 412586
rect 251804 412528 254674 412584
rect 254730 412528 254735 412584
rect 251804 412526 254735 412528
rect 254669 412523 254735 412526
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 48129 409594 48195 409597
rect 48129 409592 52164 409594
rect 48129 409536 48134 409592
rect 48190 409536 52164 409592
rect 48129 409534 52164 409536
rect 48129 409531 48195 409534
rect 254301 406738 254367 406741
rect 251804 406736 254367 406738
rect 251804 406680 254306 406736
rect 254362 406680 254367 406736
rect 251804 406678 254367 406680
rect 254301 406675 254367 406678
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 48221 403746 48287 403749
rect 48221 403744 52164 403746
rect 48221 403688 48226 403744
rect 48282 403688 52164 403744
rect 48221 403686 52164 403688
rect 48221 403683 48287 403686
rect 254485 400890 254551 400893
rect 251804 400888 254551 400890
rect 251804 400832 254490 400888
rect 254546 400832 254551 400888
rect 251804 400830 254551 400832
rect 254485 400827 254551 400830
rect 51349 397898 51415 397901
rect 51349 397896 52164 397898
rect 51349 397840 51354 397896
rect 51410 397840 52164 397896
rect 51349 397838 52164 397840
rect 51349 397835 51415 397838
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 254485 395042 254551 395045
rect 251804 395040 254551 395042
rect 251804 394984 254490 395040
rect 254546 394984 254551 395040
rect 251804 394982 254551 394984
rect 254485 394979 254551 394982
rect 48313 392050 48379 392053
rect 48313 392048 52164 392050
rect 48313 391992 48318 392048
rect 48374 391992 52164 392048
rect 48313 391990 52164 391992
rect 48313 391987 48379 391990
rect 583520 391628 584960 391868
rect 254485 389194 254551 389197
rect 251804 389192 254551 389194
rect 251804 389136 254490 389192
rect 254546 389136 254551 389192
rect 251804 389134 254551 389136
rect 254485 389131 254551 389134
rect 48313 386202 48379 386205
rect 48313 386200 52164 386202
rect 48313 386144 48318 386200
rect 48374 386144 52164 386200
rect 48313 386142 52164 386144
rect 48313 386139 48379 386142
rect -960 384284 480 384524
rect 254209 383346 254275 383349
rect 251804 383344 254275 383346
rect 251804 383288 254214 383344
rect 254270 383288 254275 383344
rect 251804 383286 254275 383288
rect 254209 383283 254275 383286
rect 49417 380354 49483 380357
rect 49417 380352 52164 380354
rect 49417 380296 49422 380352
rect 49478 380296 52164 380352
rect 49417 380294 52164 380296
rect 49417 380291 49483 380294
rect 580349 378450 580415 378453
rect 583520 378450 584960 378540
rect 580349 378448 584960 378450
rect 580349 378392 580354 378448
rect 580410 378392 584960 378448
rect 580349 378390 584960 378392
rect 580349 378387 580415 378390
rect 583520 378300 584960 378390
rect 254117 377498 254183 377501
rect 251804 377496 254183 377498
rect 251804 377440 254122 377496
rect 254178 377440 254183 377496
rect 251804 377438 254183 377440
rect 254117 377435 254183 377438
rect 48221 374506 48287 374509
rect 48221 374504 52164 374506
rect 48221 374448 48226 374504
rect 48282 374448 52164 374504
rect 48221 374446 52164 374448
rect 48221 374443 48287 374446
rect 254393 371650 254459 371653
rect 251804 371648 254459 371650
rect 251804 371592 254398 371648
rect 254454 371592 254459 371648
rect 251804 371590 254459 371592
rect 254393 371587 254459 371590
rect -960 371228 480 371468
rect 48129 368658 48195 368661
rect 48129 368656 52164 368658
rect 48129 368600 48134 368656
rect 48190 368600 52164 368656
rect 48129 368598 52164 368600
rect 48129 368595 48195 368598
rect 254485 365802 254551 365805
rect 251804 365800 254551 365802
rect 251804 365744 254490 365800
rect 254546 365744 254551 365800
rect 251804 365742 254551 365744
rect 254485 365739 254551 365742
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 48037 362810 48103 362813
rect 48037 362808 52164 362810
rect 48037 362752 48042 362808
rect 48098 362752 52164 362808
rect 48037 362750 52164 362752
rect 48037 362747 48103 362750
rect 253933 359954 253999 359957
rect 251804 359952 253999 359954
rect 251804 359896 253938 359952
rect 253994 359896 253999 359952
rect 251804 359894 253999 359896
rect 253933 359891 253999 359894
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 51349 356962 51415 356965
rect 51349 356960 52164 356962
rect 51349 356904 51354 356960
rect 51410 356904 52164 356960
rect 51349 356902 52164 356904
rect 51349 356899 51415 356902
rect 254485 354106 254551 354109
rect 251804 354104 254551 354106
rect 251804 354048 254490 354104
rect 254546 354048 254551 354104
rect 251804 354046 254551 354048
rect 254485 354043 254551 354046
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 47945 351114 48011 351117
rect 47945 351112 52164 351114
rect 47945 351056 47950 351112
rect 48006 351056 52164 351112
rect 47945 351054 52164 351056
rect 47945 351051 48011 351054
rect 254761 348258 254827 348261
rect 251804 348256 254827 348258
rect 251804 348200 254766 348256
rect 254822 348200 254827 348256
rect 251804 348198 254827 348200
rect 254761 348195 254827 348198
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 47853 345266 47919 345269
rect 47853 345264 52164 345266
rect 47853 345208 47858 345264
rect 47914 345208 52164 345264
rect 47853 345206 52164 345208
rect 47853 345203 47919 345206
rect 254669 342410 254735 342413
rect 251804 342408 254735 342410
rect 251804 342352 254674 342408
rect 254730 342352 254735 342408
rect 251804 342350 254735 342352
rect 254669 342347 254735 342350
rect 299974 340036 299980 340100
rect 300044 340098 300050 340100
rect 320909 340098 320975 340101
rect 300044 340096 320975 340098
rect 300044 340040 320914 340096
rect 320970 340040 320975 340096
rect 300044 340038 320975 340040
rect 300044 340036 300050 340038
rect 320909 340035 320975 340038
rect 51441 339418 51507 339421
rect 51441 339416 52164 339418
rect 51441 339360 51446 339416
rect 51502 339360 52164 339416
rect 51441 339358 52164 339360
rect 51441 339355 51507 339358
rect 583520 338452 584960 338692
rect 254669 336562 254735 336565
rect 251804 336560 254735 336562
rect 251804 336504 254674 336560
rect 254730 336504 254735 336560
rect 251804 336502 254735 336504
rect 254669 336499 254735 336502
rect 298502 334596 298508 334660
rect 298572 334658 298578 334660
rect 321553 334658 321619 334661
rect 298572 334656 321619 334658
rect 298572 334600 321558 334656
rect 321614 334600 321619 334656
rect 298572 334598 321619 334600
rect 298572 334596 298578 334598
rect 321553 334595 321619 334598
rect 51625 333570 51691 333573
rect 51625 333568 52164 333570
rect 51625 333512 51630 333568
rect 51686 333512 52164 333568
rect 51625 333510 52164 333512
rect 51625 333507 51691 333510
rect -960 332196 480 332436
rect 293217 332210 293283 332213
rect 310329 332210 310395 332213
rect 293217 332208 310395 332210
rect 293217 332152 293222 332208
rect 293278 332152 310334 332208
rect 310390 332152 310395 332208
rect 293217 332150 310395 332152
rect 293217 332147 293283 332150
rect 310329 332147 310395 332150
rect 253381 332074 253447 332077
rect 341885 332074 341951 332077
rect 253381 332072 341951 332074
rect 253381 332016 253386 332072
rect 253442 332016 341890 332072
rect 341946 332016 341951 332072
rect 253381 332014 341951 332016
rect 253381 332011 253447 332014
rect 341885 332011 341951 332014
rect 295926 331876 295932 331940
rect 295996 331938 296002 331940
rect 296529 331938 296595 331941
rect 295996 331936 296595 331938
rect 295996 331880 296534 331936
rect 296590 331880 296595 331936
rect 295996 331878 296595 331880
rect 295996 331876 296002 331878
rect 296529 331875 296595 331878
rect 296529 331802 296595 331805
rect 322933 331802 322999 331805
rect 296529 331800 322999 331802
rect 296529 331744 296534 331800
rect 296590 331744 322938 331800
rect 322994 331744 322999 331800
rect 296529 331742 322999 331744
rect 296529 331739 296595 331742
rect 322933 331739 322999 331742
rect 253197 331666 253263 331669
rect 300669 331666 300735 331669
rect 253197 331664 300735 331666
rect 253197 331608 253202 331664
rect 253258 331608 300674 331664
rect 300730 331608 300735 331664
rect 253197 331606 300735 331608
rect 253197 331603 253263 331606
rect 300669 331603 300735 331606
rect 293401 331530 293467 331533
rect 348969 331530 349035 331533
rect 293401 331528 349035 331530
rect 293401 331472 293406 331528
rect 293462 331472 348974 331528
rect 349030 331472 349035 331528
rect 293401 331470 349035 331472
rect 293401 331467 293467 331470
rect 348969 331467 349035 331470
rect 253565 331394 253631 331397
rect 316125 331394 316191 331397
rect 253565 331392 316191 331394
rect 253565 331336 253570 331392
rect 253626 331336 316130 331392
rect 316186 331336 316191 331392
rect 253565 331334 316191 331336
rect 253565 331331 253631 331334
rect 316125 331331 316191 331334
rect 300158 331196 300164 331260
rect 300228 331258 300234 331260
rect 305177 331258 305243 331261
rect 300228 331256 305243 331258
rect 300228 331200 305182 331256
rect 305238 331200 305243 331256
rect 300228 331198 305243 331200
rect 300228 331196 300234 331198
rect 305177 331195 305243 331198
rect 254209 330714 254275 330717
rect 251804 330712 254275 330714
rect 251804 330656 254214 330712
rect 254270 330656 254275 330712
rect 251804 330654 254275 330656
rect 254209 330651 254275 330654
rect 297357 329762 297423 329765
rect 297357 329760 300196 329762
rect 297357 329704 297362 329760
rect 297418 329704 300196 329760
rect 297357 329702 300196 329704
rect 297357 329699 297423 329702
rect 350257 329082 350323 329085
rect 349876 329080 350323 329082
rect 349876 329024 350262 329080
rect 350318 329024 350323 329080
rect 349876 329022 350323 329024
rect 350257 329019 350323 329022
rect 297449 328402 297515 328405
rect 297449 328400 300196 328402
rect 297449 328344 297454 328400
rect 297510 328344 300196 328400
rect 297449 328342 300196 328344
rect 297449 328339 297515 328342
rect 49417 327722 49483 327725
rect 350165 327722 350231 327725
rect 49417 327720 52164 327722
rect 49417 327664 49422 327720
rect 49478 327664 52164 327720
rect 49417 327662 52164 327664
rect 349876 327720 350231 327722
rect 349876 327664 350170 327720
rect 350226 327664 350231 327720
rect 349876 327662 350231 327664
rect 49417 327659 49483 327662
rect 350165 327659 350231 327662
rect 349981 326906 350047 326909
rect 349846 326904 350047 326906
rect 349846 326848 349986 326904
rect 350042 326848 350047 326904
rect 349846 326846 350047 326848
rect 297541 326362 297607 326365
rect 297541 326360 300196 326362
rect 297541 326304 297546 326360
rect 297602 326304 300196 326360
rect 349846 326332 349906 326846
rect 349981 326843 350047 326846
rect 297541 326302 300196 326304
rect 297541 326299 297607 326302
rect 580349 325274 580415 325277
rect 583520 325274 584960 325364
rect 580349 325272 584960 325274
rect 580349 325216 580354 325272
rect 580410 325216 584960 325272
rect 580349 325214 584960 325216
rect 580349 325211 580415 325214
rect 583520 325124 584960 325214
rect 297265 325002 297331 325005
rect 350073 325002 350139 325005
rect 297265 325000 300196 325002
rect 297265 324944 297270 325000
rect 297326 324944 300196 325000
rect 297265 324942 300196 324944
rect 349876 325000 350139 325002
rect 349876 324944 350078 325000
rect 350134 324944 350139 325000
rect 349876 324942 350139 324944
rect 297265 324939 297331 324942
rect 350073 324939 350139 324942
rect 254485 324866 254551 324869
rect 251804 324864 254551 324866
rect 251804 324808 254490 324864
rect 254546 324808 254551 324864
rect 251804 324806 254551 324808
rect 254485 324803 254551 324806
rect 297725 323642 297791 323645
rect 352741 323642 352807 323645
rect 297725 323640 300196 323642
rect 297725 323584 297730 323640
rect 297786 323584 300196 323640
rect 297725 323582 300196 323584
rect 349876 323640 352807 323642
rect 349876 323584 352746 323640
rect 352802 323584 352807 323640
rect 349876 323582 352807 323584
rect 297725 323579 297791 323582
rect 352741 323579 352807 323582
rect 299657 322282 299723 322285
rect 299657 322280 300196 322282
rect 299657 322224 299662 322280
rect 299718 322224 300196 322280
rect 299657 322222 300196 322224
rect 299657 322219 299723 322222
rect 49325 321874 49391 321877
rect 49325 321872 52164 321874
rect 49325 321816 49330 321872
rect 49386 321816 52164 321872
rect 49325 321814 52164 321816
rect 49325 321811 49391 321814
rect 351913 321602 351979 321605
rect 349876 321600 351979 321602
rect 349876 321544 351918 321600
rect 351974 321544 351979 321600
rect 349876 321542 351979 321544
rect 351913 321539 351979 321542
rect 297081 320242 297147 320245
rect 351862 320242 351868 320244
rect 297081 320240 300196 320242
rect 297081 320184 297086 320240
rect 297142 320184 300196 320240
rect 297081 320182 300196 320184
rect 349876 320182 351868 320242
rect 297081 320179 297147 320182
rect 351862 320180 351868 320182
rect 351932 320180 351938 320244
rect -960 319140 480 319380
rect 254301 319018 254367 319021
rect 251804 319016 254367 319018
rect 251804 318960 254306 319016
rect 254362 318960 254367 319016
rect 251804 318958 254367 318960
rect 254301 318955 254367 318958
rect 297173 318882 297239 318885
rect 352373 318882 352439 318885
rect 297173 318880 300196 318882
rect 297173 318824 297178 318880
rect 297234 318824 300196 318880
rect 297173 318822 300196 318824
rect 349876 318880 352439 318882
rect 349876 318824 352378 318880
rect 352434 318824 352439 318880
rect 349876 318822 352439 318824
rect 297173 318819 297239 318822
rect 352373 318819 352439 318822
rect 297725 317522 297791 317525
rect 350901 317522 350967 317525
rect 297725 317520 300196 317522
rect 297725 317464 297730 317520
rect 297786 317464 300196 317520
rect 297725 317462 300196 317464
rect 349876 317520 350967 317522
rect 349876 317464 350906 317520
rect 350962 317464 350967 317520
rect 349876 317462 350967 317464
rect 297725 317459 297791 317462
rect 350901 317459 350967 317462
rect 297725 316162 297791 316165
rect 297725 316160 300196 316162
rect 297725 316104 297730 316160
rect 297786 316104 300196 316160
rect 297725 316102 300196 316104
rect 297725 316099 297791 316102
rect 49233 316026 49299 316029
rect 49233 316024 52164 316026
rect 49233 315968 49238 316024
rect 49294 315968 52164 316024
rect 49233 315966 52164 315968
rect 49233 315963 49299 315966
rect 349797 315754 349863 315757
rect 349797 315752 349906 315754
rect 349797 315696 349802 315752
rect 349858 315696 349906 315752
rect 349797 315691 349906 315696
rect 349846 315452 349906 315691
rect 297909 314802 297975 314805
rect 297909 314800 300196 314802
rect 297909 314744 297914 314800
rect 297970 314744 300196 314800
rect 297909 314742 300196 314744
rect 297909 314739 297975 314742
rect 351453 314122 351519 314125
rect 349876 314120 351519 314122
rect 349876 314064 351458 314120
rect 351514 314064 351519 314120
rect 349876 314062 351519 314064
rect 351453 314059 351519 314062
rect 254669 313170 254735 313173
rect 251804 313168 254735 313170
rect 251804 313112 254674 313168
rect 254730 313112 254735 313168
rect 251804 313110 254735 313112
rect 254669 313107 254735 313110
rect 297909 312762 297975 312765
rect 297909 312760 300196 312762
rect 297909 312704 297914 312760
rect 297970 312704 300196 312760
rect 297909 312702 300196 312704
rect 297909 312699 297975 312702
rect 349846 312221 349906 312732
rect 349797 312216 349906 312221
rect 349797 312160 349802 312216
rect 349858 312160 349906 312216
rect 349797 312158 349906 312160
rect 349797 312155 349863 312158
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 298001 311402 298067 311405
rect 299238 311402 299244 311404
rect 298001 311400 299244 311402
rect 298001 311344 298006 311400
rect 298062 311344 299244 311400
rect 298001 311342 299244 311344
rect 298001 311339 298067 311342
rect 299238 311340 299244 311342
rect 299308 311402 299314 311404
rect 351913 311402 351979 311405
rect 299308 311342 300196 311402
rect 349876 311400 351979 311402
rect 349876 311344 351918 311400
rect 351974 311344 351979 311400
rect 349876 311342 351979 311344
rect 299308 311340 299314 311342
rect 351913 311339 351979 311342
rect 51533 310178 51599 310181
rect 51533 310176 52164 310178
rect 51533 310120 51538 310176
rect 51594 310120 52164 310176
rect 51533 310118 52164 310120
rect 51533 310115 51599 310118
rect 297214 309980 297220 310044
rect 297284 310042 297290 310044
rect 352373 310042 352439 310045
rect 297284 309982 300196 310042
rect 349876 310040 352439 310042
rect 349876 309984 352378 310040
rect 352434 309984 352439 310040
rect 349876 309982 352439 309984
rect 297284 309980 297290 309982
rect 352373 309979 352439 309982
rect 298645 308682 298711 308685
rect 298645 308680 300196 308682
rect 298645 308624 298650 308680
rect 298706 308624 300196 308680
rect 298645 308622 300196 308624
rect 298645 308619 298711 308622
rect 350901 308002 350967 308005
rect 349876 308000 350967 308002
rect 349876 307944 350906 308000
rect 350962 307944 350967 308000
rect 349876 307942 350967 307944
rect 350901 307939 350967 307942
rect 254209 307322 254275 307325
rect 251804 307320 254275 307322
rect 251804 307264 254214 307320
rect 254270 307264 254275 307320
rect 251804 307262 254275 307264
rect 254209 307259 254275 307262
rect 298001 306642 298067 306645
rect 352005 306642 352071 306645
rect 298001 306640 300196 306642
rect 298001 306584 298006 306640
rect 298062 306584 300196 306640
rect 298001 306582 300196 306584
rect 349876 306640 352071 306642
rect 349876 306584 352010 306640
rect 352066 306584 352071 306640
rect 349876 306582 352071 306584
rect 298001 306579 298067 306582
rect 352005 306579 352071 306582
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 349981 305826 350047 305829
rect 349846 305824 350047 305826
rect 349846 305768 349986 305824
rect 350042 305768 350047 305824
rect 349846 305766 350047 305768
rect 298001 305282 298067 305285
rect 298001 305280 300196 305282
rect 298001 305224 298006 305280
rect 298062 305224 300196 305280
rect 349846 305252 349906 305766
rect 349981 305763 350047 305766
rect 298001 305222 300196 305224
rect 298001 305219 298067 305222
rect 349889 304466 349955 304469
rect 349846 304464 349955 304466
rect 349846 304408 349894 304464
rect 349950 304408 349955 304464
rect 349846 304403 349955 304408
rect 49141 304330 49207 304333
rect 49141 304328 52164 304330
rect 49141 304272 49146 304328
rect 49202 304272 52164 304328
rect 49141 304270 52164 304272
rect 49141 304267 49207 304270
rect 298553 303922 298619 303925
rect 298553 303920 300196 303922
rect 298553 303864 298558 303920
rect 298614 303864 300196 303920
rect 349846 303892 349906 304403
rect 298553 303862 300196 303864
rect 298553 303859 298619 303862
rect 298001 302562 298067 302565
rect 298001 302560 300196 302562
rect 298001 302504 298006 302560
rect 298062 302504 300196 302560
rect 298001 302502 300196 302504
rect 298001 302499 298067 302502
rect 350717 301882 350783 301885
rect 349876 301880 350783 301882
rect 349876 301824 350722 301880
rect 350778 301824 350783 301880
rect 349876 301822 350783 301824
rect 350717 301819 350783 301822
rect 254669 301474 254735 301477
rect 251804 301472 254735 301474
rect 251804 301416 254674 301472
rect 254730 301416 254735 301472
rect 251804 301414 254735 301416
rect 254669 301411 254735 301414
rect 296989 301202 297055 301205
rect 296989 301200 300196 301202
rect 296989 301144 296994 301200
rect 297050 301144 300196 301200
rect 296989 301142 300196 301144
rect 296989 301139 297055 301142
rect 351453 300522 351519 300525
rect 349876 300520 351519 300522
rect 349876 300464 351458 300520
rect 351514 300464 351519 300520
rect 349876 300462 351519 300464
rect 351453 300459 351519 300462
rect 297817 299162 297883 299165
rect 350809 299162 350875 299165
rect 297817 299160 300196 299162
rect 297817 299104 297822 299160
rect 297878 299104 300196 299160
rect 297817 299102 300196 299104
rect 349876 299160 350875 299162
rect 349876 299104 350814 299160
rect 350870 299104 350875 299160
rect 349876 299102 350875 299104
rect 297817 299099 297883 299102
rect 350809 299099 350875 299102
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect 48681 298482 48747 298485
rect 48681 298480 52164 298482
rect 48681 298424 48686 298480
rect 48742 298424 52164 298480
rect 48681 298422 52164 298424
rect 48681 298419 48747 298422
rect 299565 297802 299631 297805
rect 352097 297802 352163 297805
rect 299565 297800 300196 297802
rect 299565 297744 299570 297800
rect 299626 297744 300196 297800
rect 299565 297742 300196 297744
rect 349876 297800 352163 297802
rect 349876 297744 352102 297800
rect 352158 297744 352163 297800
rect 349876 297742 352163 297744
rect 299565 297739 299631 297742
rect 352097 297739 352163 297742
rect 297725 296442 297791 296445
rect 352465 296442 352531 296445
rect 297725 296440 300196 296442
rect 297725 296384 297730 296440
rect 297786 296384 300196 296440
rect 297725 296382 300196 296384
rect 349876 296440 352531 296442
rect 349876 296384 352470 296440
rect 352526 296384 352531 296440
rect 349876 296382 352531 296384
rect 297725 296379 297791 296382
rect 352465 296379 352531 296382
rect 254669 295626 254735 295629
rect 251804 295624 254735 295626
rect 251804 295568 254674 295624
rect 254730 295568 254735 295624
rect 251804 295566 254735 295568
rect 254669 295563 254735 295566
rect 297817 295082 297883 295085
rect 297817 295080 300196 295082
rect 297817 295024 297822 295080
rect 297878 295024 300196 295080
rect 297817 295022 300196 295024
rect 297817 295019 297883 295022
rect 351913 294402 351979 294405
rect 349876 294400 351979 294402
rect 349876 294344 351918 294400
rect 351974 294344 351979 294400
rect 349876 294342 351979 294344
rect 351913 294339 351979 294342
rect -960 293178 480 293268
rect 3601 293178 3667 293181
rect -960 293176 3667 293178
rect -960 293120 3606 293176
rect 3662 293120 3667 293176
rect -960 293118 3667 293120
rect -960 293028 480 293118
rect 3601 293115 3667 293118
rect 352097 293042 352163 293045
rect 349876 293040 352163 293042
rect 48773 292634 48839 292637
rect 48773 292632 52164 292634
rect 48773 292576 48778 292632
rect 48834 292576 52164 292632
rect 48773 292574 52164 292576
rect 48773 292571 48839 292574
rect 284886 292572 284892 292636
rect 284956 292634 284962 292636
rect 300166 292634 300226 293012
rect 349876 292984 352102 293040
rect 352158 292984 352163 293040
rect 349876 292982 352163 292984
rect 352097 292979 352163 292982
rect 284956 292574 300226 292634
rect 284956 292572 284962 292574
rect 298001 291682 298067 291685
rect 350717 291682 350783 291685
rect 353477 291682 353543 291685
rect 298001 291680 300196 291682
rect 298001 291624 298006 291680
rect 298062 291624 300196 291680
rect 298001 291622 300196 291624
rect 349876 291680 353543 291682
rect 349876 291624 350722 291680
rect 350778 291624 353482 291680
rect 353538 291624 353543 291680
rect 349876 291622 353543 291624
rect 298001 291619 298067 291622
rect 350717 291619 350783 291622
rect 353477 291619 353543 291622
rect 297909 290322 297975 290325
rect 352281 290322 352347 290325
rect 297909 290320 300196 290322
rect 297909 290264 297914 290320
rect 297970 290264 300196 290320
rect 297909 290262 300196 290264
rect 349876 290320 352347 290322
rect 349876 290264 352286 290320
rect 352342 290264 352347 290320
rect 349876 290262 352347 290264
rect 297909 290259 297975 290262
rect 352281 290259 352347 290262
rect 254025 289778 254091 289781
rect 251804 289776 254091 289778
rect 251804 289720 254030 289776
rect 254086 289720 254091 289776
rect 251804 289718 254091 289720
rect 254025 289715 254091 289718
rect 298001 288962 298067 288965
rect 298001 288960 300196 288962
rect 298001 288904 298006 288960
rect 298062 288904 300196 288960
rect 298001 288902 300196 288904
rect 298001 288899 298067 288902
rect 351085 288282 351151 288285
rect 349876 288280 351151 288282
rect 349876 288224 351090 288280
rect 351146 288224 351151 288280
rect 349876 288222 351151 288224
rect 351085 288219 351151 288222
rect 298001 287602 298067 287605
rect 298001 287600 300196 287602
rect 298001 287544 298006 287600
rect 298062 287544 300196 287600
rect 298001 287542 300196 287544
rect 298001 287539 298067 287542
rect 351913 286922 351979 286925
rect 349876 286920 351979 286922
rect 349876 286864 351918 286920
rect 351974 286864 351979 286920
rect 349876 286862 351979 286864
rect 351913 286859 351979 286862
rect 51950 286726 52164 286786
rect 51950 286514 52010 286726
rect 52085 286514 52151 286517
rect 51950 286512 52151 286514
rect 51950 286456 52090 286512
rect 52146 286456 52151 286512
rect 51950 286454 52151 286456
rect 52085 286451 52151 286454
rect 297909 285562 297975 285565
rect 352281 285562 352347 285565
rect 297909 285560 300196 285562
rect 297909 285504 297914 285560
rect 297970 285504 300196 285560
rect 297909 285502 300196 285504
rect 349876 285560 352347 285562
rect 349876 285504 352286 285560
rect 352342 285504 352347 285560
rect 349876 285502 352347 285504
rect 297909 285499 297975 285502
rect 352281 285499 352347 285502
rect 583520 285276 584960 285516
rect 297633 284202 297699 284205
rect 350993 284202 351059 284205
rect 297633 284200 300196 284202
rect 297633 284144 297638 284200
rect 297694 284144 300196 284200
rect 297633 284142 300196 284144
rect 349876 284200 351059 284202
rect 349876 284144 350998 284200
rect 351054 284144 351059 284200
rect 349876 284142 351059 284144
rect 297633 284139 297699 284142
rect 350993 284139 351059 284142
rect 254301 283930 254367 283933
rect 251804 283928 254367 283930
rect 251804 283872 254306 283928
rect 254362 283872 254367 283928
rect 251804 283870 254367 283872
rect 254301 283867 254367 283870
rect 299565 282842 299631 282845
rect 352649 282842 352715 282845
rect 299565 282840 300196 282842
rect 299565 282784 299570 282840
rect 299626 282784 300196 282840
rect 299565 282782 300196 282784
rect 349876 282840 352715 282842
rect 349876 282784 352654 282840
rect 352710 282784 352715 282840
rect 349876 282782 352715 282784
rect 299565 282779 299631 282782
rect 352649 282779 352715 282782
rect 295425 282162 295491 282165
rect 295926 282162 295932 282164
rect 295425 282160 295932 282162
rect 295425 282104 295430 282160
rect 295486 282104 295932 282160
rect 295425 282102 295932 282104
rect 295425 282099 295491 282102
rect 295926 282100 295932 282102
rect 295996 282100 296002 282164
rect 51349 282026 51415 282029
rect 291142 282026 291148 282028
rect 51349 282024 291148 282026
rect 51349 281968 51354 282024
rect 51410 281968 291148 282024
rect 51349 281966 291148 281968
rect 51349 281963 51415 281966
rect 291142 281964 291148 281966
rect 291212 281964 291218 282028
rect 51533 281890 51599 281893
rect 285990 281890 285996 281892
rect 51533 281888 285996 281890
rect 51533 281832 51538 281888
rect 51594 281832 285996 281888
rect 51533 281830 285996 281832
rect 51533 281827 51599 281830
rect 285990 281828 285996 281830
rect 286060 281828 286066 281892
rect 299238 281420 299244 281484
rect 299308 281482 299314 281484
rect 299473 281482 299539 281485
rect 299308 281480 299539 281482
rect 299308 281424 299478 281480
rect 299534 281424 299539 281480
rect 299308 281422 299539 281424
rect 299308 281420 299314 281422
rect 299473 281419 299539 281422
rect 299614 281422 300196 281482
rect 47945 281346 48011 281349
rect 290774 281346 290780 281348
rect 47945 281344 290780 281346
rect 47945 281288 47950 281344
rect 48006 281288 290780 281344
rect 47945 281286 290780 281288
rect 47945 281283 48011 281286
rect 290774 281284 290780 281286
rect 290844 281284 290850 281348
rect 299013 281346 299079 281349
rect 299614 281346 299674 281422
rect 299013 281344 299674 281346
rect 299013 281288 299018 281344
rect 299074 281288 299674 281344
rect 299013 281286 299674 281288
rect 299013 281283 299079 281286
rect 47853 281210 47919 281213
rect 290590 281210 290596 281212
rect 47853 281208 290596 281210
rect 47853 281152 47858 281208
rect 47914 281152 290596 281208
rect 47853 281150 290596 281152
rect 47853 281147 47919 281150
rect 290590 281148 290596 281150
rect 290660 281148 290666 281212
rect 49417 281074 49483 281077
rect 287278 281074 287284 281076
rect 49417 281072 287284 281074
rect 49417 281016 49422 281072
rect 49478 281016 287284 281072
rect 49417 281014 287284 281016
rect 49417 281011 49483 281014
rect 287278 281012 287284 281014
rect 287348 281012 287354 281076
rect 49325 280938 49391 280941
rect 287462 280938 287468 280940
rect 49325 280936 287468 280938
rect 49325 280880 49330 280936
rect 49386 280880 287468 280936
rect 49325 280878 287468 280880
rect 49325 280875 49391 280878
rect 287462 280876 287468 280878
rect 287532 280876 287538 280940
rect 51441 280802 51507 280805
rect 288750 280802 288756 280804
rect 51441 280800 288756 280802
rect 51441 280744 51446 280800
rect 51502 280744 288756 280800
rect 51441 280742 288756 280744
rect 51441 280739 51507 280742
rect 288750 280740 288756 280742
rect 288820 280740 288826 280804
rect 350625 280802 350691 280805
rect 349876 280800 350691 280802
rect 349876 280744 350630 280800
rect 350686 280744 350691 280800
rect 349876 280742 350691 280744
rect 350625 280739 350691 280742
rect 51625 280666 51691 280669
rect 288382 280666 288388 280668
rect 51625 280664 288388 280666
rect 51625 280608 51630 280664
rect 51686 280608 288388 280664
rect 51625 280606 288388 280608
rect 51625 280603 51691 280606
rect 288382 280604 288388 280606
rect 288452 280604 288458 280668
rect 48129 280530 48195 280533
rect 292798 280530 292804 280532
rect 48129 280528 292804 280530
rect 48129 280472 48134 280528
rect 48190 280472 292804 280528
rect 48129 280470 292804 280472
rect 48129 280467 48195 280470
rect 292798 280468 292804 280470
rect 292868 280468 292874 280532
rect -960 279972 480 280212
rect 49366 278700 49372 278764
rect 49436 278762 49442 278764
rect 54569 278762 54635 278765
rect 49436 278760 54635 278762
rect 49436 278704 54574 278760
rect 54630 278704 54635 278760
rect 49436 278702 54635 278704
rect 49436 278700 49442 278702
rect 54569 278699 54635 278702
rect 59353 278082 59419 278085
rect 297214 278082 297220 278084
rect 59353 278080 297220 278082
rect 59353 278024 59358 278080
rect 59414 278024 297220 278080
rect 59353 278022 297220 278024
rect 59353 278019 59419 278022
rect 297214 278020 297220 278022
rect 297284 278020 297290 278084
rect 59445 276722 59511 276725
rect 351862 276722 351868 276724
rect 59445 276720 351868 276722
rect 59445 276664 59450 276720
rect 59506 276664 351868 276720
rect 59445 276662 351868 276664
rect 59445 276659 59511 276662
rect 351862 276660 351868 276662
rect 351932 276660 351938 276724
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267052 480 267292
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 49550 223484 49556 223548
rect 49620 223546 49626 223548
rect 55857 223546 55923 223549
rect 49620 223544 55923 223546
rect 49620 223488 55862 223544
rect 55918 223488 55923 223544
rect 49620 223486 55923 223488
rect 49620 223484 49626 223486
rect 55857 223483 55923 223486
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect 57830 218588 57836 218652
rect 57900 218650 57906 218652
rect 257613 218650 257679 218653
rect 57900 218648 257679 218650
rect 57900 218592 257618 218648
rect 257674 218592 257679 218648
rect 57900 218590 257679 218592
rect 57900 218588 57906 218590
rect 257613 218587 257679 218590
rect 297449 218242 297515 218245
rect 300158 218242 300164 218244
rect 297449 218240 300164 218242
rect 297449 218184 297454 218240
rect 297510 218184 300164 218240
rect 297449 218182 300164 218184
rect 297449 218179 297515 218182
rect 300158 218180 300164 218182
rect 300228 218180 300234 218244
rect 296805 217698 296871 217701
rect 296805 217696 300196 217698
rect 296805 217640 296810 217696
rect 296866 217640 300196 217696
rect 296805 217638 300196 217640
rect 296805 217635 296871 217638
rect 57053 217426 57119 217429
rect 57053 217424 60076 217426
rect 57053 217368 57058 217424
rect 57114 217368 60076 217424
rect 57053 217366 60076 217368
rect 57053 217363 57119 217366
rect 297725 216202 297791 216205
rect 297725 216200 300196 216202
rect 297725 216144 297730 216200
rect 297786 216144 300196 216200
rect 297725 216142 300196 216144
rect 297725 216139 297791 216142
rect 222837 215658 222903 215661
rect 219788 215656 222903 215658
rect 219788 215600 222842 215656
rect 222898 215600 222903 215656
rect 219788 215598 222903 215600
rect 222837 215595 222903 215598
rect -960 214828 480 215068
rect 297725 214706 297791 214709
rect 297725 214704 300196 214706
rect 297725 214648 297730 214704
rect 297786 214648 300196 214704
rect 297725 214646 300196 214648
rect 297725 214643 297791 214646
rect 60549 213890 60615 213893
rect 60549 213888 60658 213890
rect 60549 213832 60554 213888
rect 60610 213832 60658 213888
rect 60549 213827 60658 213832
rect 60598 213316 60658 213827
rect 297725 213210 297791 213213
rect 297725 213208 300196 213210
rect 297725 213152 297730 213208
rect 297786 213152 300196 213208
rect 297725 213150 300196 213152
rect 297725 213147 297791 213150
rect 222285 212802 222351 212805
rect 219788 212800 222351 212802
rect 219788 212744 222290 212800
rect 222346 212744 222351 212800
rect 219788 212742 222351 212744
rect 222285 212739 222351 212742
rect 297725 211714 297791 211717
rect 297725 211712 300196 211714
rect 297725 211656 297730 211712
rect 297786 211656 300196 211712
rect 297725 211654 300196 211656
rect 297725 211651 297791 211654
rect 297725 210218 297791 210221
rect 297725 210216 300196 210218
rect 297725 210160 297730 210216
rect 297786 210160 300196 210216
rect 297725 210158 300196 210160
rect 297725 210155 297791 210158
rect 223205 209946 223271 209949
rect 219788 209944 223271 209946
rect 219788 209888 223210 209944
rect 223266 209888 223271 209944
rect 219788 209886 223271 209888
rect 223205 209883 223271 209886
rect 57145 209266 57211 209269
rect 57145 209264 60076 209266
rect 57145 209208 57150 209264
rect 57206 209208 60076 209264
rect 57145 209206 60076 209208
rect 57145 209203 57211 209206
rect 297725 208722 297791 208725
rect 297725 208720 300196 208722
rect 297725 208664 297730 208720
rect 297786 208664 300196 208720
rect 297725 208662 300196 208664
rect 297725 208659 297791 208662
rect 297725 207226 297791 207229
rect 297725 207224 300196 207226
rect 297725 207168 297730 207224
rect 297786 207168 300196 207224
rect 297725 207166 300196 207168
rect 297725 207163 297791 207166
rect 222929 207090 222995 207093
rect 219788 207088 222995 207090
rect 219788 207032 222934 207088
rect 222990 207032 222995 207088
rect 219788 207030 222995 207032
rect 222929 207027 222995 207030
rect 297725 205730 297791 205733
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 297725 205728 300196 205730
rect 297725 205672 297730 205728
rect 297786 205672 300196 205728
rect 297725 205670 300196 205672
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 297725 205667 297791 205670
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 57329 205186 57395 205189
rect 57329 205184 60076 205186
rect 57329 205128 57334 205184
rect 57390 205128 60076 205184
rect 57329 205126 60076 205128
rect 57329 205123 57395 205126
rect 222837 204234 222903 204237
rect 219788 204232 222903 204234
rect 219788 204176 222842 204232
rect 222898 204176 222903 204232
rect 219788 204174 222903 204176
rect 222837 204171 222903 204174
rect 295977 204234 296043 204237
rect 295977 204232 300196 204234
rect 295977 204176 295982 204232
rect 296038 204176 300196 204232
rect 295977 204174 300196 204176
rect 295977 204171 296043 204174
rect 296805 202738 296871 202741
rect 296805 202736 300196 202738
rect 296805 202680 296810 202736
rect 296866 202680 300196 202736
rect 296805 202678 300196 202680
rect 296805 202675 296871 202678
rect -960 201922 480 202012
rect 3693 201922 3759 201925
rect -960 201920 3759 201922
rect -960 201864 3698 201920
rect 3754 201864 3759 201920
rect -960 201862 3759 201864
rect -960 201772 480 201862
rect 3693 201859 3759 201862
rect 223021 201378 223087 201381
rect 219788 201376 223087 201378
rect 219788 201320 223026 201376
rect 223082 201320 223087 201376
rect 219788 201318 223087 201320
rect 223021 201315 223087 201318
rect 297725 201242 297791 201245
rect 297725 201240 300196 201242
rect 297725 201184 297730 201240
rect 297786 201184 300196 201240
rect 297725 201182 300196 201184
rect 297725 201179 297791 201182
rect 57329 201106 57395 201109
rect 57329 201104 60076 201106
rect 57329 201048 57334 201104
rect 57390 201048 60076 201104
rect 57329 201046 60076 201048
rect 57329 201043 57395 201046
rect 297725 199746 297791 199749
rect 297725 199744 300196 199746
rect 297725 199688 297730 199744
rect 297786 199688 300196 199744
rect 297725 199686 300196 199688
rect 297725 199683 297791 199686
rect 222929 198522 222995 198525
rect 219788 198520 222995 198522
rect 219788 198464 222934 198520
rect 222990 198464 222995 198520
rect 219788 198462 222995 198464
rect 222929 198459 222995 198462
rect 297725 198250 297791 198253
rect 297725 198248 300196 198250
rect 297725 198192 297730 198248
rect 297786 198192 300196 198248
rect 297725 198190 300196 198192
rect 297725 198187 297791 198190
rect 57329 197026 57395 197029
rect 57329 197024 60076 197026
rect 57329 196968 57334 197024
rect 57390 196968 60076 197024
rect 57329 196966 60076 196968
rect 57329 196963 57395 196966
rect 297725 196754 297791 196757
rect 297725 196752 300196 196754
rect 297725 196696 297730 196752
rect 297786 196696 300196 196752
rect 297725 196694 300196 196696
rect 297725 196691 297791 196694
rect 223481 195666 223547 195669
rect 219788 195664 223547 195666
rect 219788 195608 223486 195664
rect 223542 195608 223547 195664
rect 219788 195606 223547 195608
rect 223481 195603 223547 195606
rect 297725 195258 297791 195261
rect 297725 195256 300196 195258
rect 297725 195200 297730 195256
rect 297786 195200 300196 195256
rect 297725 195198 300196 195200
rect 297725 195195 297791 195198
rect 297725 193762 297791 193765
rect 297725 193760 300196 193762
rect 297725 193704 297730 193760
rect 297786 193704 300196 193760
rect 297725 193702 300196 193704
rect 297725 193699 297791 193702
rect 57237 192946 57303 192949
rect 57237 192944 60076 192946
rect 57237 192888 57242 192944
rect 57298 192888 60076 192944
rect 57237 192886 60076 192888
rect 57237 192883 57303 192886
rect 223481 192810 223547 192813
rect 219788 192808 223547 192810
rect 219788 192752 223486 192808
rect 223542 192752 223547 192808
rect 219788 192750 223547 192752
rect 223481 192747 223547 192750
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 297541 192266 297607 192269
rect 297541 192264 300196 192266
rect 297541 192208 297546 192264
rect 297602 192208 300196 192264
rect 297541 192206 300196 192208
rect 297541 192203 297607 192206
rect 297725 190770 297791 190773
rect 297725 190768 300196 190770
rect 297725 190712 297730 190768
rect 297786 190712 300196 190768
rect 297725 190710 300196 190712
rect 297725 190707 297791 190710
rect 222837 189954 222903 189957
rect 219788 189952 222903 189954
rect 219788 189896 222842 189952
rect 222898 189896 222903 189952
rect 219788 189894 222903 189896
rect 222837 189891 222903 189894
rect 297541 189274 297607 189277
rect 297541 189272 300196 189274
rect 297541 189216 297546 189272
rect 297602 189216 300196 189272
rect 297541 189214 300196 189216
rect 297541 189211 297607 189214
rect -960 188866 480 188956
rect 3601 188866 3667 188869
rect -960 188864 3667 188866
rect -960 188808 3606 188864
rect 3662 188808 3667 188864
rect -960 188806 3667 188808
rect -960 188716 480 188806
rect 3601 188803 3667 188806
rect 57329 188866 57395 188869
rect 57329 188864 60076 188866
rect 57329 188808 57334 188864
rect 57390 188808 60076 188864
rect 57329 188806 60076 188808
rect 57329 188803 57395 188806
rect 297725 187778 297791 187781
rect 297725 187776 300196 187778
rect 297725 187720 297730 187776
rect 297786 187720 300196 187776
rect 297725 187718 300196 187720
rect 297725 187715 297791 187718
rect 222837 187098 222903 187101
rect 219788 187096 222903 187098
rect 219788 187040 222842 187096
rect 222898 187040 222903 187096
rect 219788 187038 222903 187040
rect 222837 187035 222903 187038
rect 297725 186282 297791 186285
rect 297725 186280 300196 186282
rect 297725 186224 297730 186280
rect 297786 186224 300196 186280
rect 297725 186222 300196 186224
rect 297725 186219 297791 186222
rect 56685 184786 56751 184789
rect 297725 184786 297791 184789
rect 56685 184784 60076 184786
rect 56685 184728 56690 184784
rect 56746 184728 60076 184784
rect 56685 184726 60076 184728
rect 297725 184784 300196 184786
rect 297725 184728 297730 184784
rect 297786 184728 300196 184784
rect 297725 184726 300196 184728
rect 56685 184723 56751 184726
rect 297725 184723 297791 184726
rect 222285 184242 222351 184245
rect 219788 184240 222351 184242
rect 219788 184184 222290 184240
rect 222346 184184 222351 184240
rect 219788 184182 222351 184184
rect 222285 184179 222351 184182
rect 297725 183290 297791 183293
rect 297725 183288 300196 183290
rect 297725 183232 297730 183288
rect 297786 183232 300196 183288
rect 297725 183230 300196 183232
rect 297725 183227 297791 183230
rect 297725 181794 297791 181797
rect 297725 181792 300196 181794
rect 297725 181736 297730 181792
rect 297786 181736 300196 181792
rect 297725 181734 300196 181736
rect 297725 181731 297791 181734
rect 223481 181386 223547 181389
rect 219788 181384 223547 181386
rect 219788 181328 223486 181384
rect 223542 181328 223547 181384
rect 219788 181326 223547 181328
rect 223481 181323 223547 181326
rect 56685 180706 56751 180709
rect 56685 180704 60076 180706
rect 56685 180648 56690 180704
rect 56746 180648 60076 180704
rect 56685 180646 60076 180648
rect 56685 180643 56751 180646
rect 297725 180298 297791 180301
rect 297725 180296 300196 180298
rect 297725 180240 297730 180296
rect 297786 180240 300196 180296
rect 297725 180238 300196 180240
rect 297725 180235 297791 180238
rect 583520 179210 584960 179300
rect 583342 179150 584960 179210
rect 583342 179074 583402 179150
rect 583520 179074 584960 179150
rect 583342 179060 584960 179074
rect 583342 179014 583586 179060
rect 297725 178802 297791 178805
rect 297725 178800 300196 178802
rect 297725 178744 297730 178800
rect 297786 178744 300196 178800
rect 297725 178742 300196 178744
rect 297725 178739 297791 178742
rect 222653 178530 222719 178533
rect 219788 178528 222719 178530
rect 219788 178472 222658 178528
rect 222714 178472 222719 178528
rect 219788 178470 222719 178472
rect 222653 178467 222719 178470
rect 355358 178060 355364 178124
rect 355428 178122 355434 178124
rect 583526 178122 583586 179014
rect 355428 178062 583586 178122
rect 355428 178060 355434 178062
rect 297725 177306 297791 177309
rect 297725 177304 300196 177306
rect 297725 177248 297730 177304
rect 297786 177248 300196 177304
rect 297725 177246 300196 177248
rect 297725 177243 297791 177246
rect 403566 177244 403572 177308
rect 403636 177306 403642 177308
rect 448605 177306 448671 177309
rect 403636 177304 448671 177306
rect 403636 177248 448610 177304
rect 448666 177248 448671 177304
rect 403636 177246 448671 177248
rect 403636 177244 403642 177246
rect 448605 177243 448671 177246
rect 57329 176626 57395 176629
rect 57329 176624 60076 176626
rect 57329 176568 57334 176624
rect 57390 176568 60076 176624
rect 57329 176566 60076 176568
rect 57329 176563 57395 176566
rect -960 175796 480 176036
rect 297725 175810 297791 175813
rect 297725 175808 300196 175810
rect 297725 175752 297730 175808
rect 297786 175752 300196 175808
rect 297725 175750 300196 175752
rect 297725 175747 297791 175750
rect 222653 175674 222719 175677
rect 219788 175672 222719 175674
rect 219788 175616 222658 175672
rect 222714 175616 222719 175672
rect 219788 175614 222719 175616
rect 222653 175611 222719 175614
rect 297725 174314 297791 174317
rect 297725 174312 300196 174314
rect 297725 174256 297730 174312
rect 297786 174256 300196 174312
rect 297725 174254 300196 174256
rect 297725 174251 297791 174254
rect 222377 172818 222443 172821
rect 219788 172816 222443 172818
rect 219788 172760 222382 172816
rect 222438 172760 222443 172816
rect 219788 172758 222443 172760
rect 222377 172755 222443 172758
rect 297725 172818 297791 172821
rect 297725 172816 300196 172818
rect 297725 172760 297730 172816
rect 297786 172760 300196 172816
rect 297725 172758 300196 172760
rect 297725 172755 297791 172758
rect 57237 172546 57303 172549
rect 57237 172544 60076 172546
rect 57237 172488 57242 172544
rect 57298 172488 60076 172544
rect 57237 172486 60076 172488
rect 57237 172483 57303 172486
rect 297725 171322 297791 171325
rect 297725 171320 300196 171322
rect 297725 171264 297730 171320
rect 297786 171264 300196 171320
rect 297725 171262 300196 171264
rect 297725 171259 297791 171262
rect 222469 169962 222535 169965
rect 219788 169960 222535 169962
rect 219788 169904 222474 169960
rect 222530 169904 222535 169960
rect 219788 169902 222535 169904
rect 222469 169899 222535 169902
rect 297725 169826 297791 169829
rect 297725 169824 300196 169826
rect 297725 169768 297730 169824
rect 297786 169768 300196 169824
rect 297725 169766 300196 169768
rect 297725 169763 297791 169766
rect 57329 168466 57395 168469
rect 57329 168464 60076 168466
rect 57329 168408 57334 168464
rect 57390 168408 60076 168464
rect 57329 168406 60076 168408
rect 57329 168403 57395 168406
rect 297725 168330 297791 168333
rect 297725 168328 300196 168330
rect 297725 168272 297730 168328
rect 297786 168272 300196 168328
rect 297725 168270 300196 168272
rect 297725 168267 297791 168270
rect 222929 167106 222995 167109
rect 219788 167104 222995 167106
rect 219788 167048 222934 167104
rect 222990 167048 222995 167104
rect 219788 167046 222995 167048
rect 222929 167043 222995 167046
rect 296805 166834 296871 166837
rect 296805 166832 300196 166834
rect 296805 166776 296810 166832
rect 296866 166776 300196 166832
rect 296805 166774 300196 166776
rect 296805 166771 296871 166774
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 297725 165338 297791 165341
rect 297725 165336 300196 165338
rect 297725 165280 297730 165336
rect 297786 165280 300196 165336
rect 297725 165278 300196 165280
rect 297725 165275 297791 165278
rect 55857 164386 55923 164389
rect 55857 164384 60076 164386
rect 55857 164328 55862 164384
rect 55918 164328 60076 164384
rect 55857 164326 60076 164328
rect 55857 164323 55923 164326
rect 223481 164250 223547 164253
rect 219788 164248 223547 164250
rect 219788 164192 223486 164248
rect 223542 164192 223547 164248
rect 219788 164190 223547 164192
rect 223481 164187 223547 164190
rect 297725 163842 297791 163845
rect 297725 163840 300196 163842
rect 297725 163784 297730 163840
rect 297786 163784 300196 163840
rect 297725 163782 300196 163784
rect 297725 163779 297791 163782
rect -960 162740 480 162980
rect 297725 162346 297791 162349
rect 297725 162344 300196 162346
rect 297725 162288 297730 162344
rect 297786 162288 300196 162344
rect 297725 162286 300196 162288
rect 297725 162283 297791 162286
rect 223021 161394 223087 161397
rect 219788 161392 223087 161394
rect 219788 161336 223026 161392
rect 223082 161336 223087 161392
rect 219788 161334 223087 161336
rect 223021 161331 223087 161334
rect 297725 160850 297791 160853
rect 297725 160848 300196 160850
rect 297725 160792 297730 160848
rect 297786 160792 300196 160848
rect 297725 160790 300196 160792
rect 297725 160787 297791 160790
rect 57053 160306 57119 160309
rect 57053 160304 60076 160306
rect 57053 160248 57058 160304
rect 57114 160248 60076 160304
rect 57053 160246 60076 160248
rect 57053 160243 57119 160246
rect 297725 159354 297791 159357
rect 297725 159352 300196 159354
rect 297725 159296 297730 159352
rect 297786 159296 300196 159352
rect 297725 159294 300196 159296
rect 297725 159291 297791 159294
rect 222929 158538 222995 158541
rect 219788 158536 222995 158538
rect 219788 158480 222934 158536
rect 222990 158480 222995 158536
rect 219788 158478 222995 158480
rect 222929 158475 222995 158478
rect 296805 157858 296871 157861
rect 296805 157856 300196 157858
rect 296805 157800 296810 157856
rect 296866 157800 300196 157856
rect 296805 157798 300196 157800
rect 296805 157795 296871 157798
rect 297725 156362 297791 156365
rect 297725 156360 300196 156362
rect 297725 156304 297730 156360
rect 297786 156304 300196 156360
rect 297725 156302 300196 156304
rect 297725 156299 297791 156302
rect 57053 156226 57119 156229
rect 57053 156224 60076 156226
rect 57053 156168 57058 156224
rect 57114 156168 60076 156224
rect 57053 156166 60076 156168
rect 57053 156163 57119 156166
rect 223481 155682 223547 155685
rect 219788 155680 223547 155682
rect 219788 155624 223486 155680
rect 223542 155624 223547 155680
rect 219788 155622 223547 155624
rect 223481 155619 223547 155622
rect 297725 154866 297791 154869
rect 297725 154864 300196 154866
rect 297725 154808 297730 154864
rect 297786 154808 300196 154864
rect 297725 154806 300196 154808
rect 297725 154803 297791 154806
rect 297725 153370 297791 153373
rect 297725 153368 300196 153370
rect 297725 153312 297730 153368
rect 297786 153312 300196 153368
rect 297725 153310 300196 153312
rect 297725 153307 297791 153310
rect 222561 152826 222627 152829
rect 219788 152824 222627 152826
rect 219788 152768 222566 152824
rect 222622 152768 222627 152824
rect 219788 152766 222627 152768
rect 222561 152763 222627 152766
rect 579797 152690 579863 152693
rect 583520 152690 584960 152780
rect 579797 152688 584960 152690
rect 579797 152632 579802 152688
rect 579858 152632 584960 152688
rect 579797 152630 584960 152632
rect 579797 152627 579863 152630
rect 583520 152540 584960 152630
rect 57329 152146 57395 152149
rect 57329 152144 60076 152146
rect 57329 152088 57334 152144
rect 57390 152088 60076 152144
rect 57329 152086 60076 152088
rect 57329 152083 57395 152086
rect 297725 151874 297791 151877
rect 297725 151872 300196 151874
rect 297725 151816 297730 151872
rect 297786 151816 300196 151872
rect 297725 151814 300196 151816
rect 297725 151811 297791 151814
rect 297725 150378 297791 150381
rect 297725 150376 300196 150378
rect 297725 150320 297730 150376
rect 297786 150320 300196 150376
rect 297725 150318 300196 150320
rect 297725 150315 297791 150318
rect 223481 149970 223547 149973
rect 219788 149968 223547 149970
rect -960 149834 480 149924
rect 219788 149912 223486 149968
rect 223542 149912 223547 149968
rect 219788 149910 223547 149912
rect 223481 149907 223547 149910
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 296805 148882 296871 148885
rect 296805 148880 300196 148882
rect 296805 148824 296810 148880
rect 296866 148824 300196 148880
rect 296805 148822 300196 148824
rect 296805 148819 296871 148822
rect 57329 148066 57395 148069
rect 57329 148064 60076 148066
rect 57329 148008 57334 148064
rect 57390 148008 60076 148064
rect 57329 148006 60076 148008
rect 57329 148003 57395 148006
rect 341057 147522 341123 147525
rect 339940 147520 341123 147522
rect 339940 147464 341062 147520
rect 341118 147464 341123 147520
rect 339940 147462 341123 147464
rect 341057 147459 341123 147462
rect 297725 147386 297791 147389
rect 297725 147384 300196 147386
rect 297725 147328 297730 147384
rect 297786 147328 300196 147384
rect 297725 147326 300196 147328
rect 297725 147323 297791 147326
rect 223481 147114 223547 147117
rect 219788 147112 223547 147114
rect 219788 147056 223486 147112
rect 223542 147056 223547 147112
rect 219788 147054 223547 147056
rect 223481 147051 223547 147054
rect 297725 145890 297791 145893
rect 297725 145888 300196 145890
rect 297725 145832 297730 145888
rect 297786 145832 300196 145888
rect 297725 145830 300196 145832
rect 297725 145827 297791 145830
rect 340137 145346 340203 145349
rect 339940 145344 340203 145346
rect 339940 145288 340142 145344
rect 340198 145288 340203 145344
rect 339940 145286 340203 145288
rect 340137 145283 340203 145286
rect 297725 144394 297791 144397
rect 297725 144392 300196 144394
rect 297725 144336 297730 144392
rect 297786 144336 300196 144392
rect 297725 144334 300196 144336
rect 297725 144331 297791 144334
rect 222469 144258 222535 144261
rect 219788 144256 222535 144258
rect 219788 144200 222474 144256
rect 222530 144200 222535 144256
rect 219788 144198 222535 144200
rect 222469 144195 222535 144198
rect 57329 143986 57395 143989
rect 57329 143984 60076 143986
rect 57329 143928 57334 143984
rect 57390 143928 60076 143984
rect 57329 143926 60076 143928
rect 57329 143923 57395 143926
rect 342253 143170 342319 143173
rect 339940 143168 342319 143170
rect 339940 143112 342258 143168
rect 342314 143112 342319 143168
rect 339940 143110 342319 143112
rect 342253 143107 342319 143110
rect 297541 142898 297607 142901
rect 297541 142896 300196 142898
rect 297541 142840 297546 142896
rect 297602 142840 300196 142896
rect 297541 142838 300196 142840
rect 297541 142835 297607 142838
rect 223481 141402 223547 141405
rect 219788 141400 223547 141402
rect 219788 141344 223486 141400
rect 223542 141344 223547 141400
rect 219788 141342 223547 141344
rect 223481 141339 223547 141342
rect 297725 141402 297791 141405
rect 297725 141400 300196 141402
rect 297725 141344 297730 141400
rect 297786 141344 300196 141400
rect 297725 141342 300196 141344
rect 297725 141339 297791 141342
rect 340873 140994 340939 140997
rect 339940 140992 340939 140994
rect 339940 140936 340878 140992
rect 340934 140936 340939 140992
rect 339940 140934 340939 140936
rect 340873 140931 340939 140934
rect 57421 139906 57487 139909
rect 297725 139906 297791 139909
rect 57421 139904 60076 139906
rect 57421 139848 57426 139904
rect 57482 139848 60076 139904
rect 57421 139846 60076 139848
rect 297725 139904 300196 139906
rect 297725 139848 297730 139904
rect 297786 139848 300196 139904
rect 297725 139846 300196 139848
rect 57421 139843 57487 139846
rect 297725 139843 297791 139846
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 339940 138758 340154 138818
rect 340094 138685 340154 138758
rect 340045 138680 340154 138685
rect 340045 138624 340050 138680
rect 340106 138624 340154 138680
rect 340045 138622 340154 138624
rect 340045 138619 340111 138622
rect 222929 138546 222995 138549
rect 219788 138544 222995 138546
rect 219788 138488 222934 138544
rect 222990 138488 222995 138544
rect 219788 138486 222995 138488
rect 222929 138483 222995 138486
rect 297725 138410 297791 138413
rect 297725 138408 300196 138410
rect 297725 138352 297730 138408
rect 297786 138352 300196 138408
rect 297725 138350 300196 138352
rect 297725 138347 297791 138350
rect 297725 136914 297791 136917
rect 297725 136912 300196 136914
rect -960 136778 480 136868
rect 297725 136856 297730 136912
rect 297786 136856 300196 136912
rect 297725 136854 300196 136856
rect 297725 136851 297791 136854
rect 3141 136778 3207 136781
rect -960 136776 3207 136778
rect -960 136720 3146 136776
rect 3202 136720 3207 136776
rect -960 136718 3207 136720
rect -960 136628 480 136718
rect 3141 136715 3207 136718
rect 342345 136642 342411 136645
rect 339940 136640 342411 136642
rect 339940 136584 342350 136640
rect 342406 136584 342411 136640
rect 339940 136582 342411 136584
rect 342345 136579 342411 136582
rect 57329 135826 57395 135829
rect 57329 135824 60076 135826
rect 57329 135768 57334 135824
rect 57390 135768 60076 135824
rect 57329 135766 60076 135768
rect 57329 135763 57395 135766
rect 222837 135690 222903 135693
rect 219788 135688 222903 135690
rect 219788 135632 222842 135688
rect 222898 135632 222903 135688
rect 219788 135630 222903 135632
rect 222837 135627 222903 135630
rect 296805 135418 296871 135421
rect 296805 135416 300196 135418
rect 296805 135360 296810 135416
rect 296866 135360 300196 135416
rect 296805 135358 300196 135360
rect 296805 135355 296871 135358
rect 342437 134466 342503 134469
rect 339940 134464 342503 134466
rect 339940 134408 342442 134464
rect 342498 134408 342503 134464
rect 339940 134406 342503 134408
rect 342437 134403 342503 134406
rect 297725 133922 297791 133925
rect 297725 133920 300196 133922
rect 297725 133864 297730 133920
rect 297786 133864 300196 133920
rect 297725 133862 300196 133864
rect 297725 133859 297791 133862
rect 222469 132834 222535 132837
rect 219788 132832 222535 132834
rect 219788 132776 222474 132832
rect 222530 132776 222535 132832
rect 219788 132774 222535 132776
rect 222469 132771 222535 132774
rect 297725 132426 297791 132429
rect 297725 132424 300196 132426
rect 297725 132368 297730 132424
rect 297786 132368 300196 132424
rect 297725 132366 300196 132368
rect 297725 132363 297791 132366
rect 341241 132290 341307 132293
rect 339940 132288 341307 132290
rect 339940 132232 341246 132288
rect 341302 132232 341307 132288
rect 339940 132230 341307 132232
rect 341241 132227 341307 132230
rect 57830 131684 57836 131748
rect 57900 131746 57906 131748
rect 57900 131686 60076 131746
rect 57900 131684 57906 131686
rect 297725 130930 297791 130933
rect 297725 130928 300196 130930
rect 297725 130872 297730 130928
rect 297786 130872 300196 130928
rect 297725 130870 300196 130872
rect 297725 130867 297791 130870
rect 342529 130114 342595 130117
rect 339940 130112 342595 130114
rect 339940 130056 342534 130112
rect 342590 130056 342595 130112
rect 339940 130054 342595 130056
rect 342529 130051 342595 130054
rect 223113 129978 223179 129981
rect 219788 129976 223179 129978
rect 219788 129920 223118 129976
rect 223174 129920 223179 129976
rect 219788 129918 223179 129920
rect 223113 129915 223179 129918
rect 297725 129434 297791 129437
rect 297725 129432 300196 129434
rect 297725 129376 297730 129432
rect 297786 129376 300196 129432
rect 297725 129374 300196 129376
rect 297725 129371 297791 129374
rect 297725 127938 297791 127941
rect 342621 127938 342687 127941
rect 297725 127936 300196 127938
rect 297725 127880 297730 127936
rect 297786 127880 300196 127936
rect 297725 127878 300196 127880
rect 339940 127936 342687 127938
rect 339940 127880 342626 127936
rect 342682 127880 342687 127936
rect 339940 127878 342687 127880
rect 297725 127875 297791 127878
rect 342621 127875 342687 127878
rect 58893 127666 58959 127669
rect 58893 127664 60076 127666
rect 58893 127608 58898 127664
rect 58954 127608 60076 127664
rect 58893 127606 60076 127608
rect 58893 127603 58959 127606
rect 223481 127122 223547 127125
rect 219788 127120 223547 127122
rect 219788 127064 223486 127120
rect 223542 127064 223547 127120
rect 219788 127062 223547 127064
rect 223481 127059 223547 127062
rect 297725 126442 297791 126445
rect 297725 126440 300196 126442
rect 297725 126384 297730 126440
rect 297786 126384 300196 126440
rect 297725 126382 300196 126384
rect 297725 126379 297791 126382
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 342713 125762 342779 125765
rect 339940 125760 342779 125762
rect 339940 125704 342718 125760
rect 342774 125704 342779 125760
rect 339940 125702 342779 125704
rect 342713 125699 342779 125702
rect 297725 124946 297791 124949
rect 297725 124944 300196 124946
rect 297725 124888 297730 124944
rect 297786 124888 300196 124944
rect 297725 124886 300196 124888
rect 297725 124883 297791 124886
rect 222469 124266 222535 124269
rect 219788 124264 222535 124266
rect 219788 124208 222474 124264
rect 222530 124208 222535 124264
rect 219788 124206 222535 124208
rect 222469 124203 222535 124206
rect -960 123572 480 123812
rect 57513 123586 57579 123589
rect 342805 123586 342871 123589
rect 57513 123584 60076 123586
rect 57513 123528 57518 123584
rect 57574 123528 60076 123584
rect 57513 123526 60076 123528
rect 339940 123584 342871 123586
rect 339940 123528 342810 123584
rect 342866 123528 342871 123584
rect 339940 123526 342871 123528
rect 57513 123523 57579 123526
rect 342805 123523 342871 123526
rect 297725 123450 297791 123453
rect 297725 123448 300196 123450
rect 297725 123392 297730 123448
rect 297786 123392 300196 123448
rect 297725 123390 300196 123392
rect 297725 123387 297791 123390
rect 297725 121954 297791 121957
rect 297725 121952 300196 121954
rect 297725 121896 297730 121952
rect 297786 121896 300196 121952
rect 297725 121894 300196 121896
rect 297725 121891 297791 121894
rect 223205 121410 223271 121413
rect 341149 121410 341215 121413
rect 219788 121408 223271 121410
rect 219788 121352 223210 121408
rect 223266 121352 223271 121408
rect 219788 121350 223271 121352
rect 339940 121408 341215 121410
rect 339940 121352 341154 121408
rect 341210 121352 341215 121408
rect 339940 121350 341215 121352
rect 223205 121347 223271 121350
rect 341149 121347 341215 121350
rect 297725 120458 297791 120461
rect 297725 120456 300196 120458
rect 297725 120400 297730 120456
rect 297786 120400 300196 120456
rect 297725 120398 300196 120400
rect 297725 120395 297791 120398
rect 58801 119506 58867 119509
rect 58801 119504 60076 119506
rect 58801 119448 58806 119504
rect 58862 119448 60076 119504
rect 58801 119446 60076 119448
rect 58801 119443 58867 119446
rect 340229 119234 340295 119237
rect 339940 119232 340295 119234
rect 339940 119176 340234 119232
rect 340290 119176 340295 119232
rect 339940 119174 340295 119176
rect 340229 119171 340295 119174
rect 297725 118962 297791 118965
rect 297725 118960 300196 118962
rect 297725 118904 297730 118960
rect 297786 118904 300196 118960
rect 297725 118902 300196 118904
rect 297725 118899 297791 118902
rect 223481 118554 223547 118557
rect 219788 118552 223547 118554
rect 219788 118496 223486 118552
rect 223542 118496 223547 118552
rect 219788 118494 223547 118496
rect 223481 118491 223547 118494
rect 296805 117466 296871 117469
rect 296805 117464 300196 117466
rect 296805 117408 296810 117464
rect 296866 117408 300196 117464
rect 296805 117406 300196 117408
rect 296805 117403 296871 117406
rect 342897 117058 342963 117061
rect 339940 117056 342963 117058
rect 339940 117000 342902 117056
rect 342958 117000 342963 117056
rect 339940 116998 342963 117000
rect 342897 116995 342963 116998
rect 297725 115970 297791 115973
rect 297725 115968 300196 115970
rect 297725 115912 297730 115968
rect 297786 115912 300196 115968
rect 297725 115910 300196 115912
rect 297725 115907 297791 115910
rect 223481 115698 223547 115701
rect 219788 115696 223547 115698
rect 219788 115640 223486 115696
rect 223542 115640 223547 115696
rect 219788 115638 223547 115640
rect 223481 115635 223547 115638
rect 59537 115426 59603 115429
rect 59537 115424 60076 115426
rect 59537 115368 59542 115424
rect 59598 115368 60076 115424
rect 59537 115366 60076 115368
rect 59537 115363 59603 115366
rect 340965 114882 341031 114885
rect 339940 114880 341031 114882
rect 339940 114824 340970 114880
rect 341026 114824 341031 114880
rect 339940 114822 341031 114824
rect 340965 114819 341031 114822
rect 297725 114474 297791 114477
rect 297725 114472 300196 114474
rect 297725 114416 297730 114472
rect 297786 114416 300196 114472
rect 297725 114414 300196 114416
rect 297725 114411 297791 114414
rect 297725 112978 297791 112981
rect 297725 112976 300196 112978
rect 297725 112920 297730 112976
rect 297786 112920 300196 112976
rect 297725 112918 300196 112920
rect 297725 112915 297791 112918
rect 222193 112842 222259 112845
rect 219788 112840 222259 112842
rect 219788 112784 222198 112840
rect 222254 112784 222259 112840
rect 219788 112782 222259 112784
rect 222193 112779 222259 112782
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 341333 112706 341399 112709
rect 339940 112704 341399 112706
rect 339940 112648 341338 112704
rect 341394 112648 341399 112704
rect 583520 112692 584960 112782
rect 339940 112646 341399 112648
rect 341333 112643 341399 112646
rect 299105 111482 299171 111485
rect 299105 111480 300196 111482
rect 299105 111424 299110 111480
rect 299166 111424 300196 111480
rect 299105 111422 300196 111424
rect 299105 111419 299171 111422
rect 58985 111346 59051 111349
rect 58985 111344 60076 111346
rect 58985 111288 58990 111344
rect 59046 111288 60076 111344
rect 58985 111286 60076 111288
rect 58985 111283 59051 111286
rect -960 110516 480 110756
rect 340321 110530 340387 110533
rect 339940 110528 340387 110530
rect 339940 110472 340326 110528
rect 340382 110472 340387 110528
rect 339940 110470 340387 110472
rect 340321 110467 340387 110470
rect 223481 109986 223547 109989
rect 219788 109984 223547 109986
rect 219788 109928 223486 109984
rect 223542 109928 223547 109984
rect 219788 109926 223547 109928
rect 223481 109923 223547 109926
rect 297265 109986 297331 109989
rect 297265 109984 300196 109986
rect 297265 109928 297270 109984
rect 297326 109928 300196 109984
rect 297265 109926 300196 109928
rect 297265 109923 297331 109926
rect 299197 108490 299263 108493
rect 299197 108488 300196 108490
rect 299197 108432 299202 108488
rect 299258 108432 300196 108488
rect 299197 108430 300196 108432
rect 299197 108427 299263 108430
rect 340822 108354 340828 108356
rect 339940 108294 340828 108354
rect 340822 108292 340828 108294
rect 340892 108354 340898 108356
rect 342897 108354 342963 108357
rect 340892 108352 342963 108354
rect 340892 108296 342902 108352
rect 342958 108296 342963 108352
rect 340892 108294 342963 108296
rect 340892 108292 340898 108294
rect 342897 108291 342963 108294
rect 57605 107266 57671 107269
rect 57605 107264 60076 107266
rect 57605 107208 57610 107264
rect 57666 107208 60076 107264
rect 57605 107206 60076 107208
rect 57605 107203 57671 107206
rect 222653 107130 222719 107133
rect 219788 107128 222719 107130
rect 219788 107072 222658 107128
rect 222714 107072 222719 107128
rect 219788 107070 222719 107072
rect 222653 107067 222719 107070
rect 297909 106994 297975 106997
rect 297909 106992 300196 106994
rect 297909 106936 297914 106992
rect 297970 106936 300196 106992
rect 297909 106934 300196 106936
rect 297909 106931 297975 106934
rect 342294 106178 342300 106180
rect 339940 106118 342300 106178
rect 342294 106116 342300 106118
rect 342364 106178 342370 106180
rect 342897 106178 342963 106181
rect 342364 106176 342963 106178
rect 342364 106120 342902 106176
rect 342958 106120 342963 106176
rect 342364 106118 342963 106120
rect 342364 106116 342370 106118
rect 342897 106115 342963 106118
rect 299289 105498 299355 105501
rect 299289 105496 300196 105498
rect 299289 105440 299294 105496
rect 299350 105440 300196 105496
rect 299289 105438 300196 105440
rect 299289 105435 299355 105438
rect 222837 104274 222903 104277
rect 219788 104272 222903 104274
rect 219788 104216 222842 104272
rect 222898 104216 222903 104272
rect 219788 104214 222903 104216
rect 222837 104211 222903 104214
rect 297357 104002 297423 104005
rect 341425 104002 341491 104005
rect 297357 104000 300196 104002
rect 297357 103944 297362 104000
rect 297418 103944 300196 104000
rect 297357 103942 300196 103944
rect 339940 104000 341491 104002
rect 339940 103944 341430 104000
rect 341486 103944 341491 104000
rect 339940 103942 341491 103944
rect 297357 103939 297423 103942
rect 341425 103939 341491 103942
rect 57697 103186 57763 103189
rect 57697 103184 60076 103186
rect 57697 103128 57702 103184
rect 57758 103128 60076 103184
rect 57697 103126 60076 103128
rect 57697 103123 57763 103126
rect 296989 102506 297055 102509
rect 296989 102504 300196 102506
rect 296989 102448 296994 102504
rect 297050 102448 300196 102504
rect 296989 102446 300196 102448
rect 296989 102443 297055 102446
rect 341517 101826 341583 101829
rect 339940 101824 341583 101826
rect 339940 101768 341522 101824
rect 341578 101768 341583 101824
rect 339940 101766 341583 101768
rect 341517 101763 341583 101766
rect 223481 101418 223547 101421
rect 219788 101416 223547 101418
rect 219788 101360 223486 101416
rect 223542 101360 223547 101416
rect 219788 101358 223547 101360
rect 223481 101355 223547 101358
rect 297633 101010 297699 101013
rect 297633 101008 300196 101010
rect 297633 100952 297638 101008
rect 297694 100952 300196 101008
rect 297633 100950 300196 100952
rect 297633 100947 297699 100950
rect 341609 99650 341675 99653
rect 339940 99648 341675 99650
rect 339940 99592 341614 99648
rect 341670 99592 341675 99648
rect 339940 99590 341675 99592
rect 341609 99587 341675 99590
rect 297449 99514 297515 99517
rect 580257 99514 580323 99517
rect 583520 99514 584960 99604
rect 297449 99512 300196 99514
rect 297449 99456 297454 99512
rect 297510 99456 300196 99512
rect 297449 99454 300196 99456
rect 580257 99512 584960 99514
rect 580257 99456 580262 99512
rect 580318 99456 584960 99512
rect 580257 99454 584960 99456
rect 297449 99451 297515 99454
rect 580257 99451 580323 99454
rect 583520 99364 584960 99454
rect 59813 99106 59879 99109
rect 59813 99104 60076 99106
rect 59813 99048 59818 99104
rect 59874 99048 60076 99104
rect 59813 99046 60076 99048
rect 59813 99043 59879 99046
rect 223021 98562 223087 98565
rect 219788 98560 223087 98562
rect 219788 98504 223026 98560
rect 223082 98504 223087 98560
rect 219788 98502 223087 98504
rect 223021 98499 223087 98502
rect 298829 98018 298895 98021
rect 298829 98016 300196 98018
rect 298829 97960 298834 98016
rect 298890 97960 300196 98016
rect 298829 97958 300196 97960
rect 298829 97955 298895 97958
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 341701 97474 341767 97477
rect 339940 97472 341767 97474
rect 339940 97416 341706 97472
rect 341762 97416 341767 97472
rect 339940 97414 341767 97416
rect 341701 97411 341767 97414
rect 297817 96522 297883 96525
rect 297817 96520 300196 96522
rect 297817 96464 297822 96520
rect 297878 96464 300196 96520
rect 297817 96462 300196 96464
rect 297817 96459 297883 96462
rect 223113 95706 223179 95709
rect 219788 95704 223179 95706
rect 219788 95648 223118 95704
rect 223174 95648 223179 95704
rect 219788 95646 223179 95648
rect 223113 95643 223179 95646
rect 341006 95298 341012 95300
rect 339940 95238 341012 95298
rect 341006 95236 341012 95238
rect 341076 95236 341082 95300
rect 59445 95026 59511 95029
rect 299381 95026 299447 95029
rect 59445 95024 60076 95026
rect 59445 94968 59450 95024
rect 59506 94968 60076 95024
rect 59445 94966 60076 94968
rect 299381 95024 300196 95026
rect 299381 94968 299386 95024
rect 299442 94968 300196 95024
rect 299381 94966 300196 94968
rect 59445 94963 59511 94966
rect 299381 94963 299447 94966
rect 298921 93530 298987 93533
rect 298921 93528 300196 93530
rect 298921 93472 298926 93528
rect 298982 93472 300196 93528
rect 298921 93470 300196 93472
rect 298921 93467 298987 93470
rect 343081 93122 343147 93125
rect 339940 93120 343147 93122
rect 339940 93064 343086 93120
rect 343142 93064 343147 93120
rect 339940 93062 343147 93064
rect 343081 93059 343147 93062
rect 223481 92850 223547 92853
rect 219788 92848 223547 92850
rect 219788 92792 223486 92848
rect 223542 92792 223547 92848
rect 219788 92790 223547 92792
rect 223481 92787 223547 92790
rect 297081 92034 297147 92037
rect 297081 92032 300196 92034
rect 297081 91976 297086 92032
rect 297142 91976 300196 92032
rect 297081 91974 300196 91976
rect 297081 91971 297147 91974
rect 59261 90946 59327 90949
rect 343173 90946 343239 90949
rect 59261 90944 60076 90946
rect 59261 90888 59266 90944
rect 59322 90888 60076 90944
rect 59261 90886 60076 90888
rect 339940 90944 343239 90946
rect 339940 90888 343178 90944
rect 343234 90888 343239 90944
rect 339940 90886 343239 90888
rect 59261 90883 59327 90886
rect 343173 90883 343239 90886
rect 298001 90538 298067 90541
rect 298001 90536 300196 90538
rect 298001 90480 298006 90536
rect 298062 90480 300196 90536
rect 298001 90478 300196 90480
rect 298001 90475 298067 90478
rect 223481 89994 223547 89997
rect 219788 89992 223547 89994
rect 219788 89936 223486 89992
rect 223542 89936 223547 89992
rect 219788 89934 223547 89936
rect 223481 89931 223547 89934
rect 299013 89042 299079 89045
rect 299013 89040 300196 89042
rect 299013 88984 299018 89040
rect 299074 88984 300196 89040
rect 299013 88982 300196 88984
rect 299013 88979 299079 88982
rect 342989 88770 343055 88773
rect 339940 88768 343055 88770
rect 339940 88712 342994 88768
rect 343050 88712 343055 88768
rect 339940 88710 343055 88712
rect 342989 88707 343055 88710
rect 298001 87546 298067 87549
rect 298001 87544 300196 87546
rect 298001 87488 298006 87544
rect 298062 87488 300196 87544
rect 298001 87486 300196 87488
rect 298001 87483 298067 87486
rect 223389 87138 223455 87141
rect 219788 87136 223455 87138
rect 219788 87080 223394 87136
rect 223450 87080 223455 87136
rect 219788 87078 223455 87080
rect 223389 87075 223455 87078
rect 57789 86866 57855 86869
rect 57789 86864 60076 86866
rect 57789 86808 57794 86864
rect 57850 86808 60076 86864
rect 57789 86806 60076 86808
rect 57789 86803 57855 86806
rect 342897 86594 342963 86597
rect 339940 86592 342963 86594
rect 339940 86536 342902 86592
rect 342958 86536 342963 86592
rect 339940 86534 342963 86536
rect 342897 86531 342963 86534
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 296805 86050 296871 86053
rect 296805 86048 300196 86050
rect 296805 85992 296810 86048
rect 296866 85992 300196 86048
rect 583520 86036 584960 86126
rect 296805 85990 300196 85992
rect 296805 85987 296871 85990
rect 340086 85444 340092 85508
rect 340156 85506 340162 85508
rect 342294 85506 342300 85508
rect 340156 85446 342300 85506
rect 340156 85444 340162 85446
rect 342294 85444 342300 85446
rect 342364 85444 342370 85508
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 297541 84554 297607 84557
rect 297541 84552 300196 84554
rect 297541 84496 297546 84552
rect 297602 84496 300196 84552
rect 297541 84494 300196 84496
rect 297541 84491 297607 84494
rect 342478 84418 342484 84420
rect 339940 84358 342484 84418
rect 342478 84356 342484 84358
rect 342548 84356 342554 84420
rect 223481 84282 223547 84285
rect 219788 84280 223547 84282
rect 219788 84224 223486 84280
rect 223542 84224 223547 84280
rect 219788 84222 223547 84224
rect 223481 84219 223547 84222
rect 297909 83058 297975 83061
rect 297909 83056 300196 83058
rect 297909 83000 297914 83056
rect 297970 83000 300196 83056
rect 297909 82998 300196 83000
rect 297909 82995 297975 82998
rect 59077 82786 59143 82789
rect 59077 82784 60076 82786
rect 59077 82728 59082 82784
rect 59138 82728 60076 82784
rect 59077 82726 60076 82728
rect 59077 82723 59143 82726
rect 342294 82242 342300 82244
rect 339940 82182 342300 82242
rect 342294 82180 342300 82182
rect 342364 82180 342370 82244
rect 297909 81562 297975 81565
rect 297909 81560 300196 81562
rect 297909 81504 297914 81560
rect 297970 81504 300196 81560
rect 297909 81502 300196 81504
rect 297909 81499 297975 81502
rect 223481 81426 223547 81429
rect 219788 81424 223547 81426
rect 219788 81368 223486 81424
rect 223542 81368 223547 81424
rect 219788 81366 223547 81368
rect 223481 81363 223547 81366
rect 298001 80066 298067 80069
rect 342529 80066 342595 80069
rect 298001 80064 300196 80066
rect 298001 80008 298006 80064
rect 298062 80008 300196 80064
rect 298001 80006 300196 80008
rect 339940 80064 342595 80066
rect 339940 80008 342534 80064
rect 342590 80008 342595 80064
rect 339940 80006 342595 80008
rect 298001 80003 298067 80006
rect 342529 80003 342595 80006
rect 341374 79324 341380 79388
rect 341444 79386 341450 79388
rect 343081 79386 343147 79389
rect 341444 79384 343147 79386
rect 341444 79328 343086 79384
rect 343142 79328 343147 79384
rect 341444 79326 343147 79328
rect 341444 79324 341450 79326
rect 343081 79323 343147 79326
rect 57881 78706 57947 78709
rect 57881 78704 60076 78706
rect 57881 78648 57886 78704
rect 57942 78648 60076 78704
rect 57881 78646 60076 78648
rect 57881 78643 57947 78646
rect 222469 78570 222535 78573
rect 219788 78568 222535 78570
rect 219788 78512 222474 78568
rect 222530 78512 222535 78568
rect 219788 78510 222535 78512
rect 222469 78507 222535 78510
rect 297541 78570 297607 78573
rect 297541 78568 300196 78570
rect 297541 78512 297546 78568
rect 297602 78512 300196 78568
rect 297541 78510 300196 78512
rect 297541 78507 297607 78510
rect 342662 77890 342668 77892
rect 339940 77830 342668 77890
rect 342662 77828 342668 77830
rect 342732 77828 342738 77892
rect 297173 77074 297239 77077
rect 297173 77072 300196 77074
rect 297173 77016 297178 77072
rect 297234 77016 300196 77072
rect 297173 77014 300196 77016
rect 297173 77011 297239 77014
rect 222193 75714 222259 75717
rect 340505 75714 340571 75717
rect 219788 75712 222259 75714
rect 219788 75656 222198 75712
rect 222254 75656 222259 75712
rect 219788 75654 222259 75656
rect 339940 75712 340571 75714
rect 339940 75656 340510 75712
rect 340566 75656 340571 75712
rect 339940 75654 340571 75656
rect 222193 75651 222259 75654
rect 340505 75651 340571 75654
rect 298001 75578 298067 75581
rect 298001 75576 300196 75578
rect 298001 75520 298006 75576
rect 298062 75520 300196 75576
rect 298001 75518 300196 75520
rect 298001 75515 298067 75518
rect 59721 74626 59787 74629
rect 59721 74624 60076 74626
rect 59721 74568 59726 74624
rect 59782 74568 60076 74624
rect 59721 74566 60076 74568
rect 59721 74563 59787 74566
rect 298001 74082 298067 74085
rect 298001 74080 300196 74082
rect 298001 74024 298006 74080
rect 298062 74024 300196 74080
rect 298001 74022 300196 74024
rect 298001 74019 298067 74022
rect 340086 73538 340092 73540
rect 339940 73478 340092 73538
rect 340086 73476 340092 73478
rect 340156 73476 340162 73540
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 222193 72858 222259 72861
rect 219788 72856 222259 72858
rect 219788 72800 222198 72856
rect 222254 72800 222259 72856
rect 583520 72844 584960 72934
rect 219788 72798 222259 72800
rect 222193 72795 222259 72798
rect 296805 72586 296871 72589
rect 296805 72584 300196 72586
rect 296805 72528 296810 72584
rect 296866 72528 300196 72584
rect 296805 72526 300196 72528
rect 296805 72523 296871 72526
rect -960 71484 480 71724
rect 341190 71362 341196 71364
rect 339940 71302 341196 71362
rect 341190 71300 341196 71302
rect 341260 71300 341266 71364
rect 279366 71028 279372 71092
rect 279436 71090 279442 71092
rect 279436 71030 300196 71090
rect 279436 71028 279442 71030
rect 59353 70546 59419 70549
rect 59353 70544 60076 70546
rect 59353 70488 59358 70544
rect 59414 70488 60076 70544
rect 59353 70486 60076 70488
rect 59353 70483 59419 70486
rect 223481 70002 223547 70005
rect 219788 70000 223547 70002
rect 219788 69944 223486 70000
rect 223542 69944 223547 70000
rect 219788 69942 223547 69944
rect 223481 69939 223547 69942
rect 298001 69594 298067 69597
rect 298001 69592 300196 69594
rect 298001 69536 298006 69592
rect 298062 69536 300196 69592
rect 298001 69534 300196 69536
rect 298001 69531 298067 69534
rect 343081 69186 343147 69189
rect 339940 69184 343147 69186
rect 339940 69128 343086 69184
rect 343142 69128 343147 69184
rect 339940 69126 343147 69128
rect 343081 69123 343147 69126
rect 297173 68098 297239 68101
rect 297173 68096 300196 68098
rect 297173 68040 297178 68096
rect 297234 68040 300196 68096
rect 297173 68038 300196 68040
rect 297173 68035 297239 68038
rect 223481 67146 223547 67149
rect 219788 67144 223547 67146
rect 219788 67088 223486 67144
rect 223542 67088 223547 67144
rect 219788 67086 223547 67088
rect 223481 67083 223547 67086
rect 343173 67010 343239 67013
rect 339940 67008 343239 67010
rect 339940 66952 343178 67008
rect 343234 66952 343239 67008
rect 339940 66950 343239 66952
rect 343173 66947 343239 66950
rect 297541 66602 297607 66605
rect 297541 66600 300196 66602
rect 297541 66544 297546 66600
rect 297602 66544 300196 66600
rect 297541 66542 300196 66544
rect 297541 66539 297607 66542
rect 59629 66466 59695 66469
rect 59629 66464 60076 66466
rect 59629 66408 59634 66464
rect 59690 66408 60076 66464
rect 59629 66406 60076 66408
rect 59629 66403 59695 66406
rect 297357 65106 297423 65109
rect 297357 65104 300196 65106
rect 297357 65048 297362 65104
rect 297418 65048 300196 65104
rect 297357 65046 300196 65048
rect 297357 65043 297423 65046
rect 343173 64834 343239 64837
rect 339940 64832 343239 64834
rect 339940 64776 343178 64832
rect 343234 64776 343239 64832
rect 339940 64774 343239 64776
rect 343173 64771 343239 64774
rect 222837 64290 222903 64293
rect 219788 64288 222903 64290
rect 219788 64232 222842 64288
rect 222898 64232 222903 64288
rect 219788 64230 222903 64232
rect 222837 64227 222903 64230
rect 297909 63610 297975 63613
rect 297909 63608 300196 63610
rect 297909 63552 297914 63608
rect 297970 63552 300196 63608
rect 297909 63550 300196 63552
rect 297909 63547 297975 63550
rect 342345 62658 342411 62661
rect 339940 62656 342411 62658
rect 339940 62600 342350 62656
rect 342406 62600 342411 62656
rect 339940 62598 342411 62600
rect 342345 62595 342411 62598
rect 59169 62386 59235 62389
rect 59169 62384 60076 62386
rect 59169 62328 59174 62384
rect 59230 62328 60076 62384
rect 59169 62326 60076 62328
rect 59169 62323 59235 62326
rect 298001 62114 298067 62117
rect 298001 62112 300196 62114
rect 298001 62056 298006 62112
rect 298062 62056 300196 62112
rect 298001 62054 300196 62056
rect 298001 62051 298067 62054
rect 126973 61434 127039 61437
rect 341190 61434 341196 61436
rect 126973 61432 341196 61434
rect 126973 61376 126978 61432
rect 127034 61376 341196 61432
rect 126973 61374 341196 61376
rect 126973 61371 127039 61374
rect 341190 61372 341196 61374
rect 341260 61372 341266 61436
rect 317413 60346 317479 60349
rect 349654 60346 349660 60348
rect 317413 60344 349660 60346
rect 317413 60288 317418 60344
rect 317474 60288 349660 60344
rect 317413 60286 349660 60288
rect 317413 60283 317479 60286
rect 349654 60284 349660 60286
rect 349724 60284 349730 60348
rect 165613 60210 165679 60213
rect 341006 60210 341012 60212
rect 165613 60208 341012 60210
rect 165613 60152 165618 60208
rect 165674 60152 341012 60208
rect 165613 60150 341012 60152
rect 165613 60147 165679 60150
rect 341006 60148 341012 60150
rect 341076 60148 341082 60212
rect 136633 60074 136699 60077
rect 342662 60074 342668 60076
rect 136633 60072 342668 60074
rect 136633 60016 136638 60072
rect 136694 60016 342668 60072
rect 136633 60014 342668 60016
rect 136633 60011 136699 60014
rect 342662 60012 342668 60014
rect 342732 60012 342738 60076
rect 129733 59938 129799 59941
rect 339534 59938 339540 59940
rect 129733 59936 339540 59938
rect 129733 59880 129738 59936
rect 129794 59880 339540 59936
rect 129733 59878 339540 59880
rect 129733 59875 129799 59878
rect 339534 59876 339540 59878
rect 339604 59876 339610 59940
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 147673 58578 147739 58581
rect 342478 58578 342484 58580
rect 147673 58576 342484 58578
rect 147673 58520 147678 58576
rect 147734 58520 342484 58576
rect 147673 58518 342484 58520
rect 147673 58515 147739 58518
rect 342478 58516 342484 58518
rect 342548 58516 342554 58580
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 489678 39204 489684 39268
rect 489748 39266 489754 39268
rect 495433 39266 495499 39269
rect 489748 39264 495499 39266
rect 489748 39208 495438 39264
rect 495494 39208 495499 39264
rect 489748 39206 495499 39208
rect 489748 39204 489754 39206
rect 495433 39203 495499 39206
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 355174 19348 355180 19412
rect 355244 19410 355250 19412
rect 583526 19410 583586 19622
rect 355244 19350 583586 19410
rect 355244 19348 355250 19350
rect 143533 10434 143599 10437
rect 342294 10434 342300 10436
rect 143533 10432 342300 10434
rect 143533 10376 143538 10432
rect 143594 10376 342300 10432
rect 143533 10374 342300 10376
rect 143533 10371 143599 10374
rect 342294 10372 342300 10374
rect 342364 10372 342370 10436
rect 95785 10298 95851 10301
rect 508998 10298 509004 10300
rect 95785 10296 509004 10298
rect 95785 10240 95790 10296
rect 95846 10240 509004 10296
rect 95785 10238 509004 10240
rect 95785 10235 95851 10238
rect 508998 10236 509004 10238
rect 509068 10236 509074 10300
rect 74993 8938 75059 8941
rect 503662 8938 503668 8940
rect 74993 8936 503668 8938
rect 74993 8880 74998 8936
rect 75054 8880 503668 8936
rect 74993 8878 503668 8880
rect 74993 8875 75059 8878
rect 503662 8876 503668 8878
rect 503732 8876 503738 8940
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 4061 6490 4127 6493
rect -960 6488 4127 6490
rect -960 6432 4066 6488
rect 4122 6432 4127 6488
rect 583520 6476 584960 6566
rect -960 6430 4127 6432
rect -960 6340 480 6430
rect 4061 6427 4127 6430
rect 187325 4858 187391 4861
rect 340822 4858 340828 4860
rect 187325 4856 340828 4858
rect 187325 4800 187330 4856
rect 187386 4800 340828 4856
rect 187325 4798 340828 4800
rect 187325 4795 187391 4798
rect 340822 4796 340828 4798
rect 340892 4796 340898 4860
rect 484158 3980 484164 4044
rect 484228 4042 484234 4044
rect 492305 4042 492371 4045
rect 484228 4040 492371 4042
rect 484228 3984 492310 4040
rect 492366 3984 492371 4040
rect 484228 3982 492371 3984
rect 484228 3980 484234 3982
rect 492305 3979 492371 3982
rect 297265 3634 297331 3637
rect 298502 3634 298508 3636
rect 297265 3632 298508 3634
rect 297265 3576 297270 3632
rect 297326 3576 298508 3632
rect 297265 3574 298508 3576
rect 297265 3571 297331 3574
rect 298502 3572 298508 3574
rect 298572 3572 298578 3636
rect 299974 3572 299980 3636
rect 300044 3634 300050 3636
rect 300761 3634 300827 3637
rect 300044 3632 300827 3634
rect 300044 3576 300766 3632
rect 300822 3576 300827 3632
rect 300044 3574 300827 3576
rect 300044 3572 300050 3574
rect 300761 3571 300827 3574
rect 329189 3634 329255 3637
rect 349102 3634 349108 3636
rect 329189 3632 349108 3634
rect 329189 3576 329194 3632
rect 329250 3576 349108 3632
rect 329189 3574 349108 3576
rect 329189 3571 329255 3574
rect 349102 3572 349108 3574
rect 349172 3572 349178 3636
rect 183737 3498 183803 3501
rect 340086 3498 340092 3500
rect 183737 3496 340092 3498
rect 183737 3440 183742 3496
rect 183798 3440 340092 3496
rect 183737 3438 340092 3440
rect 183737 3435 183803 3438
rect 340086 3436 340092 3438
rect 340156 3436 340162 3500
rect 162485 3362 162551 3365
rect 341374 3362 341380 3364
rect 162485 3360 341380 3362
rect 162485 3304 162490 3360
rect 162546 3304 341380 3360
rect 162485 3302 341380 3304
rect 162485 3299 162551 3302
rect 341374 3300 341380 3302
rect 341444 3300 341450 3364
<< via3 >>
rect 279372 670652 279436 670716
rect 283420 663172 283484 663236
rect 286180 663036 286244 663100
rect 317644 662900 317708 662964
rect 403020 662764 403084 662828
rect 481588 662628 481652 662692
rect 495388 662492 495452 662556
rect 290964 661812 291028 661876
rect 295932 661676 295996 661740
rect 304212 661540 304276 661604
rect 305500 661404 305564 661468
rect 49372 661268 49436 661332
rect 308628 661268 308692 661332
rect 401548 661328 401612 661332
rect 401548 661272 401598 661328
rect 401598 661272 401612 661328
rect 401548 661268 401612 661272
rect 49556 661132 49620 661196
rect 309364 661132 309428 661196
rect 512132 661132 512196 661196
rect 309180 660996 309244 661060
rect 484900 660996 484964 661060
rect 499436 660996 499500 661060
rect 291700 660588 291764 660652
rect 295012 660452 295076 660516
rect 299980 660316 300044 660380
rect 308812 660180 308876 660244
rect 489132 660180 489196 660244
rect 49188 660044 49252 660108
rect 310468 660044 310532 660108
rect 311940 659908 312004 659972
rect 50108 659832 50172 659836
rect 50108 659776 50158 659832
rect 50158 659776 50172 659832
rect 50108 659772 50172 659776
rect 297220 659772 297284 659836
rect 502012 659772 502076 659836
rect 49740 659696 49804 659700
rect 49740 659640 49790 659696
rect 49790 659640 49804 659696
rect 49740 659636 49804 659640
rect 49924 659636 49988 659700
rect 51212 659696 51276 659700
rect 51212 659640 51262 659696
rect 51262 659640 51276 659696
rect 51212 659636 51276 659640
rect 359412 642092 359476 642156
rect 398604 641956 398668 642020
rect 293172 641820 293236 641884
rect 311020 641684 311084 641748
rect 363460 641684 363524 641748
rect 307524 640868 307588 640932
rect 355364 640460 355428 640524
rect 355180 640324 355244 640388
rect 303476 639508 303540 639572
rect 362540 639916 362604 639980
rect 362356 639508 362420 639572
rect 298324 639372 298388 639436
rect 362724 639372 362788 639436
rect 364012 639432 364076 639436
rect 364012 639376 364062 639432
rect 364062 639376 364076 639432
rect 364012 639372 364076 639376
rect 282684 639236 282748 639300
rect 285444 639296 285508 639300
rect 285444 639240 285458 639296
rect 285458 639240 285508 639296
rect 285444 639236 285508 639240
rect 288204 639296 288268 639300
rect 288204 639240 288254 639296
rect 288254 639240 288268 639296
rect 288204 639236 288268 639240
rect 289492 639236 289556 639300
rect 298508 639296 298572 639300
rect 298508 639240 298522 639296
rect 298522 639240 298572 639296
rect 298508 639236 298572 639240
rect 302004 638964 302068 639028
rect 50108 618292 50172 618356
rect 49188 614212 49252 614276
rect 49188 612716 49252 612780
rect 49372 608364 49436 608428
rect 49372 607140 49436 607204
rect 49924 605916 49988 605980
rect 49556 602516 49620 602580
rect 49556 600748 49620 600812
rect 302004 600672 302068 600676
rect 302004 600616 302018 600672
rect 302018 600616 302068 600672
rect 302004 600612 302068 600616
rect 303476 600672 303540 600676
rect 303476 600616 303490 600672
rect 303490 600616 303540 600672
rect 303476 600612 303540 600616
rect 307524 600672 307588 600676
rect 307524 600616 307574 600672
rect 307574 600616 307588 600672
rect 307524 600612 307588 600616
rect 360700 598300 360764 598364
rect 366220 598164 366284 598228
rect 369900 598164 369964 598228
rect 379284 598164 379348 598228
rect 373212 597620 373276 597684
rect 362540 596804 362604 596868
rect 404860 596804 404924 596868
rect 382780 595444 382844 595508
rect 373396 592588 373460 592652
rect 392532 586332 392596 586396
rect 364012 585652 364076 585716
rect 387012 583748 387076 583812
rect 362540 583068 362604 583132
rect 388300 582932 388364 582996
rect 391980 581844 392044 581908
rect 368244 581708 368308 581772
rect 380940 581572 381004 581636
rect 371740 580348 371804 580412
rect 376156 580212 376220 580276
rect 282684 578988 282748 579052
rect 311020 578852 311084 578916
rect 384068 576812 384132 576876
rect 391060 574772 391124 574836
rect 389588 574636 389652 574700
rect 396580 573276 396644 573340
rect 370084 571916 370148 571980
rect 362356 569196 362420 569260
rect 376892 568108 376956 568172
rect 368428 567972 368492 568036
rect 376340 567972 376404 568036
rect 279372 567836 279436 567900
rect 380572 566340 380636 566404
rect 49740 565796 49804 565860
rect 361620 565116 361684 565180
rect 373764 564980 373828 565044
rect 279372 564572 279436 564636
rect 361436 563892 361500 563956
rect 400260 563756 400324 563820
rect 285444 563620 285508 563684
rect 398788 563620 398852 563684
rect 298324 562260 298388 562324
rect 399156 562260 399220 562324
rect 362724 561036 362788 561100
rect 364748 560900 364812 560964
rect 362908 560220 362972 560284
rect 385540 560220 385604 560284
rect 298508 559540 298572 559604
rect 363460 558860 363524 558924
rect 400444 558180 400508 558244
rect 401732 555324 401796 555388
rect 359044 554236 359108 554300
rect 289492 554100 289556 554164
rect 400628 554100 400692 554164
rect 358860 553964 358924 554028
rect 358308 553420 358372 553484
rect 403572 552060 403636 552124
rect 358676 551924 358740 551988
rect 358492 551788 358556 551852
rect 293172 551516 293236 551580
rect 288204 551380 288268 551444
rect 400812 551380 400876 551444
rect 398972 551244 399036 551308
rect 358124 550564 358188 550628
rect 399340 550564 399404 550628
rect 401548 549204 401612 549268
rect 400812 547708 400876 547772
rect 358308 547028 358372 547092
rect 399340 543764 399404 543828
rect 317644 543628 317708 543692
rect 290964 543356 291028 543420
rect 295932 543220 295996 543284
rect 286180 543084 286244 543148
rect 283420 542948 283484 543012
rect 291700 542812 291764 542876
rect 311940 542812 312004 542876
rect 308628 542676 308692 542740
rect 295012 542540 295076 542604
rect 305500 542540 305564 542604
rect 309364 542540 309428 542604
rect 297220 542464 297284 542468
rect 297220 542408 297234 542464
rect 297234 542408 297284 542464
rect 297220 542404 297284 542408
rect 299980 542464 300044 542468
rect 299980 542408 299994 542464
rect 299994 542408 300044 542464
rect 299980 542404 300044 542408
rect 304212 542404 304276 542468
rect 308812 542404 308876 542468
rect 309180 542404 309244 542468
rect 310468 542404 310532 542468
rect 359044 541044 359108 541108
rect 358124 540636 358188 540700
rect 287284 539684 287348 539748
rect 49188 539548 49252 539612
rect 284892 539548 284956 539612
rect 285996 539548 286060 539612
rect 287468 539548 287532 539612
rect 288388 539548 288452 539612
rect 288756 539548 288820 539612
rect 290596 539608 290660 539612
rect 290596 539552 290610 539608
rect 290610 539552 290660 539608
rect 290596 539548 290660 539552
rect 290780 539608 290844 539612
rect 290780 539552 290830 539608
rect 290830 539552 290844 539608
rect 290780 539548 290844 539552
rect 291148 539548 291212 539612
rect 292804 539548 292868 539612
rect 403020 539548 403084 539612
rect 400628 537780 400692 537844
rect 399340 535604 399404 535668
rect 399340 533156 399404 533220
rect 481588 532612 481652 532676
rect 484900 532612 484964 532676
rect 489132 532612 489196 532676
rect 502012 532612 502076 532676
rect 499436 532476 499500 532540
rect 358492 530572 358556 530636
rect 484164 529892 484228 529956
rect 489684 529484 489748 529548
rect 502380 529544 502444 529548
rect 502380 529488 502430 529544
rect 502430 529488 502444 529544
rect 502380 529484 502444 529488
rect 503668 529484 503732 529548
rect 509372 527444 509436 527508
rect 360516 526900 360580 526964
rect 49372 521656 49436 521660
rect 49372 521600 49386 521656
rect 49386 521600 49436 521656
rect 49372 521596 49436 521600
rect 399340 521596 399404 521660
rect 349108 518876 349172 518940
rect 399340 518740 399404 518804
rect 512132 512756 512196 512820
rect 404860 509416 404924 509420
rect 404860 509360 404910 509416
rect 404910 509360 404924 509416
rect 404860 509356 404924 509360
rect 401732 508268 401796 508332
rect 399340 507724 399404 507788
rect 358860 505004 358924 505068
rect 400444 504800 400508 504864
rect 49556 503100 49620 503164
rect 358676 502284 358740 502348
rect 400260 501400 400324 501464
rect 359412 501196 359476 501260
rect 361436 499836 361500 499900
rect 361620 499836 361684 499900
rect 364748 499836 364812 499900
rect 368244 499836 368308 499900
rect 368612 499836 368676 499900
rect 370084 499836 370148 499900
rect 373764 499836 373828 499900
rect 376340 499836 376404 499900
rect 376892 499836 376956 499900
rect 380572 499896 380636 499900
rect 380572 499840 380622 499896
rect 380622 499840 380636 499896
rect 380572 499836 380636 499840
rect 380940 499836 381004 499900
rect 382780 499836 382844 499900
rect 385540 499836 385604 499900
rect 389588 499836 389652 499900
rect 391980 499836 392044 499900
rect 396580 499836 396644 499900
rect 392532 499700 392596 499764
rect 398604 499700 398668 499764
rect 495388 499836 495452 499900
rect 391060 499564 391124 499628
rect 366220 499428 366284 499492
rect 373212 499428 373276 499492
rect 376156 499428 376220 499492
rect 302004 499156 302068 499220
rect 369900 498884 369964 498948
rect 502380 498748 502444 498812
rect 349660 498204 349724 498268
rect 362540 498068 362604 498132
rect 384068 498068 384132 498132
rect 388300 498068 388364 498132
rect 371740 497932 371804 497996
rect 379284 497932 379348 497996
rect 362908 497796 362972 497860
rect 387012 497660 387076 497724
rect 373396 497252 373460 497316
rect 49556 484332 49620 484396
rect 51212 479708 51276 479772
rect 49372 477532 49436 477596
rect 51212 477532 51276 477596
rect 299980 340036 300044 340100
rect 298508 334596 298572 334660
rect 295932 331876 295996 331940
rect 300164 331196 300228 331260
rect 351868 320180 351932 320244
rect 299244 311340 299308 311404
rect 297220 309980 297284 310044
rect 284892 292572 284956 292636
rect 295932 282100 295996 282164
rect 291148 281964 291212 282028
rect 285996 281828 286060 281892
rect 299244 281420 299308 281484
rect 290780 281284 290844 281348
rect 290596 281148 290660 281212
rect 287284 281012 287348 281076
rect 287468 280876 287532 280940
rect 288756 280740 288820 280804
rect 288388 280604 288452 280668
rect 292804 280468 292868 280532
rect 49372 278700 49436 278764
rect 297220 278020 297284 278084
rect 351868 276660 351932 276724
rect 49556 223484 49620 223548
rect 57836 218588 57900 218652
rect 300164 218180 300228 218244
rect 355364 178060 355428 178124
rect 403572 177244 403636 177308
rect 57836 131684 57900 131748
rect 340828 108292 340892 108356
rect 342300 106116 342364 106180
rect 341012 95236 341076 95300
rect 340092 85444 340156 85508
rect 342300 85444 342364 85508
rect 342484 84356 342548 84420
rect 342300 82180 342364 82244
rect 341380 79324 341444 79388
rect 342668 77828 342732 77892
rect 340092 73476 340156 73540
rect 341196 71300 341260 71364
rect 279372 71028 279436 71092
rect 341196 61372 341260 61436
rect 349660 60284 349724 60348
rect 341012 60148 341076 60212
rect 342668 60012 342732 60076
rect 339540 59876 339604 59940
rect 342484 58516 342548 58580
rect 489684 39204 489748 39268
rect 355180 19348 355244 19412
rect 342300 10372 342364 10436
rect 509004 10236 509068 10300
rect 503668 8876 503732 8940
rect 340828 4796 340892 4860
rect 484164 3980 484228 4044
rect 298508 3572 298572 3636
rect 299980 3572 300044 3636
rect 349108 3572 349172 3636
rect 340092 3436 340156 3500
rect 341380 3300 341444 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 664000 51914 664398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 664000 56414 668898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 664000 60914 673398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 664000 65414 677898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 664000 69914 682398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 664000 74414 686898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 664000 78914 691398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 664000 83414 695898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 664000 87914 664398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 664000 92414 668898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 664000 96914 673398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 664000 101414 677898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 664000 105914 682398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 664000 110414 686898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 664000 114914 691398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 664000 119414 695898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 664000 123914 664398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 664000 128414 668898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 664000 132914 673398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 664000 137414 677898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 664000 141914 682398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 664000 146414 686898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 664000 150914 691398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 664000 155414 695898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 664000 159914 664398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 664000 164414 668898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 664000 168914 673398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 664000 173414 677898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 664000 177914 682398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 664000 182414 686898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 664000 186914 691398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 664000 191414 695898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 664000 195914 664398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 664000 200414 668898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 664000 204914 673398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 664000 209414 677898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 664000 213914 682398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 664000 218414 686898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 664000 222914 691398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 664000 227414 695898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 664000 231914 664398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 664000 236414 668898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 664000 240914 673398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 664000 245414 677898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 664000 249914 682398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 664000 254414 686898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 49371 661332 49437 661333
rect 49371 661268 49372 661332
rect 49436 661268 49437 661332
rect 49371 661267 49437 661268
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 49187 660108 49253 660109
rect 49187 660044 49188 660108
rect 49252 660044 49253 660108
rect 49187 660043 49253 660044
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 49190 614277 49250 660043
rect 49187 614276 49253 614277
rect 49187 614212 49188 614276
rect 49252 614212 49253 614276
rect 49187 614211 49253 614212
rect 49187 612780 49253 612781
rect 49187 612716 49188 612780
rect 49252 612716 49253 612780
rect 49187 612715 49253 612716
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 49190 539613 49250 612715
rect 49374 608429 49434 661267
rect 49555 661196 49621 661197
rect 49555 661132 49556 661196
rect 49620 661132 49621 661196
rect 49555 661131 49621 661132
rect 49371 608428 49437 608429
rect 49371 608364 49372 608428
rect 49436 608364 49437 608428
rect 49371 608363 49437 608364
rect 49371 607204 49437 607205
rect 49371 607140 49372 607204
rect 49436 607140 49437 607204
rect 49371 607139 49437 607140
rect 49187 539612 49253 539613
rect 49187 539548 49188 539612
rect 49252 539548 49253 539612
rect 49187 539547 49253 539548
rect 49374 521661 49434 607139
rect 49558 602581 49618 661131
rect 50107 659836 50173 659837
rect 50107 659772 50108 659836
rect 50172 659772 50173 659836
rect 50107 659771 50173 659772
rect 49739 659700 49805 659701
rect 49739 659636 49740 659700
rect 49804 659636 49805 659700
rect 49739 659635 49805 659636
rect 49923 659700 49989 659701
rect 49923 659636 49924 659700
rect 49988 659636 49989 659700
rect 49923 659635 49989 659636
rect 49555 602580 49621 602581
rect 49555 602516 49556 602580
rect 49620 602516 49621 602580
rect 49555 602515 49621 602516
rect 49555 600812 49621 600813
rect 49555 600748 49556 600812
rect 49620 600748 49621 600812
rect 49555 600747 49621 600748
rect 49371 521660 49437 521661
rect 49371 521596 49372 521660
rect 49436 521596 49437 521660
rect 49371 521595 49437 521596
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 49558 503165 49618 600747
rect 49742 565861 49802 659635
rect 49926 605981 49986 659635
rect 50110 618357 50170 659771
rect 51211 659700 51277 659701
rect 51211 659636 51212 659700
rect 51276 659636 51277 659700
rect 51211 659635 51277 659636
rect 50107 618356 50173 618357
rect 50107 618292 50108 618356
rect 50172 618292 50173 618356
rect 50107 618291 50173 618292
rect 49923 605980 49989 605981
rect 49923 605916 49924 605980
rect 49988 605916 49989 605980
rect 49923 605915 49989 605916
rect 49739 565860 49805 565861
rect 49739 565796 49740 565860
rect 49804 565796 49805 565860
rect 49739 565795 49805 565796
rect 49555 503164 49621 503165
rect 49555 503100 49556 503164
rect 49620 503100 49621 503164
rect 49555 503099 49621 503100
rect 49555 484396 49621 484397
rect 49555 484332 49556 484396
rect 49620 484332 49621 484396
rect 49555 484331 49621 484332
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 49371 477596 49437 477597
rect 49371 477532 49372 477596
rect 49436 477532 49437 477596
rect 49371 477531 49437 477532
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 49374 278765 49434 477531
rect 49371 278764 49437 278765
rect 49371 278700 49372 278764
rect 49436 278700 49437 278764
rect 49371 278699 49437 278700
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 49558 223549 49618 484331
rect 51214 479773 51274 659635
rect 71568 655954 71888 655986
rect 71568 655718 71610 655954
rect 71846 655718 71888 655954
rect 71568 655634 71888 655718
rect 71568 655398 71610 655634
rect 71846 655398 71888 655634
rect 71568 655366 71888 655398
rect 102288 655954 102608 655986
rect 102288 655718 102330 655954
rect 102566 655718 102608 655954
rect 102288 655634 102608 655718
rect 102288 655398 102330 655634
rect 102566 655398 102608 655634
rect 102288 655366 102608 655398
rect 133008 655954 133328 655986
rect 133008 655718 133050 655954
rect 133286 655718 133328 655954
rect 133008 655634 133328 655718
rect 133008 655398 133050 655634
rect 133286 655398 133328 655634
rect 133008 655366 133328 655398
rect 163728 655954 164048 655986
rect 163728 655718 163770 655954
rect 164006 655718 164048 655954
rect 163728 655634 164048 655718
rect 163728 655398 163770 655634
rect 164006 655398 164048 655634
rect 163728 655366 164048 655398
rect 194448 655954 194768 655986
rect 194448 655718 194490 655954
rect 194726 655718 194768 655954
rect 194448 655634 194768 655718
rect 194448 655398 194490 655634
rect 194726 655398 194768 655634
rect 194448 655366 194768 655398
rect 225168 655954 225488 655986
rect 225168 655718 225210 655954
rect 225446 655718 225488 655954
rect 225168 655634 225488 655718
rect 225168 655398 225210 655634
rect 225446 655398 225488 655634
rect 225168 655366 225488 655398
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 56208 651454 56528 651486
rect 56208 651218 56250 651454
rect 56486 651218 56528 651454
rect 56208 651134 56528 651218
rect 56208 650898 56250 651134
rect 56486 650898 56528 651134
rect 56208 650866 56528 650898
rect 86928 651454 87248 651486
rect 86928 651218 86970 651454
rect 87206 651218 87248 651454
rect 86928 651134 87248 651218
rect 86928 650898 86970 651134
rect 87206 650898 87248 651134
rect 86928 650866 87248 650898
rect 117648 651454 117968 651486
rect 117648 651218 117690 651454
rect 117926 651218 117968 651454
rect 117648 651134 117968 651218
rect 117648 650898 117690 651134
rect 117926 650898 117968 651134
rect 117648 650866 117968 650898
rect 148368 651454 148688 651486
rect 148368 651218 148410 651454
rect 148646 651218 148688 651454
rect 148368 651134 148688 651218
rect 148368 650898 148410 651134
rect 148646 650898 148688 651134
rect 148368 650866 148688 650898
rect 179088 651454 179408 651486
rect 179088 651218 179130 651454
rect 179366 651218 179408 651454
rect 179088 651134 179408 651218
rect 179088 650898 179130 651134
rect 179366 650898 179408 651134
rect 179088 650866 179408 650898
rect 209808 651454 210128 651486
rect 209808 651218 209850 651454
rect 210086 651218 210128 651454
rect 209808 651134 210128 651218
rect 209808 650898 209850 651134
rect 210086 650898 210128 651134
rect 209808 650866 210128 650898
rect 240528 651454 240848 651486
rect 240528 651218 240570 651454
rect 240806 651218 240848 651454
rect 240528 651134 240848 651218
rect 240528 650898 240570 651134
rect 240806 650898 240848 651134
rect 240528 650866 240848 650898
rect 71568 619954 71888 619986
rect 71568 619718 71610 619954
rect 71846 619718 71888 619954
rect 71568 619634 71888 619718
rect 71568 619398 71610 619634
rect 71846 619398 71888 619634
rect 71568 619366 71888 619398
rect 102288 619954 102608 619986
rect 102288 619718 102330 619954
rect 102566 619718 102608 619954
rect 102288 619634 102608 619718
rect 102288 619398 102330 619634
rect 102566 619398 102608 619634
rect 102288 619366 102608 619398
rect 133008 619954 133328 619986
rect 133008 619718 133050 619954
rect 133286 619718 133328 619954
rect 133008 619634 133328 619718
rect 133008 619398 133050 619634
rect 133286 619398 133328 619634
rect 133008 619366 133328 619398
rect 163728 619954 164048 619986
rect 163728 619718 163770 619954
rect 164006 619718 164048 619954
rect 163728 619634 164048 619718
rect 163728 619398 163770 619634
rect 164006 619398 164048 619634
rect 163728 619366 164048 619398
rect 194448 619954 194768 619986
rect 194448 619718 194490 619954
rect 194726 619718 194768 619954
rect 194448 619634 194768 619718
rect 194448 619398 194490 619634
rect 194726 619398 194768 619634
rect 194448 619366 194768 619398
rect 225168 619954 225488 619986
rect 225168 619718 225210 619954
rect 225446 619718 225488 619954
rect 225168 619634 225488 619718
rect 225168 619398 225210 619634
rect 225446 619398 225488 619634
rect 225168 619366 225488 619398
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 56208 615454 56528 615486
rect 56208 615218 56250 615454
rect 56486 615218 56528 615454
rect 56208 615134 56528 615218
rect 56208 614898 56250 615134
rect 56486 614898 56528 615134
rect 56208 614866 56528 614898
rect 86928 615454 87248 615486
rect 86928 615218 86970 615454
rect 87206 615218 87248 615454
rect 86928 615134 87248 615218
rect 86928 614898 86970 615134
rect 87206 614898 87248 615134
rect 86928 614866 87248 614898
rect 117648 615454 117968 615486
rect 117648 615218 117690 615454
rect 117926 615218 117968 615454
rect 117648 615134 117968 615218
rect 117648 614898 117690 615134
rect 117926 614898 117968 615134
rect 117648 614866 117968 614898
rect 148368 615454 148688 615486
rect 148368 615218 148410 615454
rect 148646 615218 148688 615454
rect 148368 615134 148688 615218
rect 148368 614898 148410 615134
rect 148646 614898 148688 615134
rect 148368 614866 148688 614898
rect 179088 615454 179408 615486
rect 179088 615218 179130 615454
rect 179366 615218 179408 615454
rect 179088 615134 179408 615218
rect 179088 614898 179130 615134
rect 179366 614898 179408 615134
rect 179088 614866 179408 614898
rect 209808 615454 210128 615486
rect 209808 615218 209850 615454
rect 210086 615218 210128 615454
rect 209808 615134 210128 615218
rect 209808 614898 209850 615134
rect 210086 614898 210128 615134
rect 209808 614866 210128 614898
rect 240528 615454 240848 615486
rect 240528 615218 240570 615454
rect 240806 615218 240848 615454
rect 240528 615134 240848 615218
rect 240528 614898 240570 615134
rect 240806 614898 240848 615134
rect 240528 614866 240848 614898
rect 71568 583954 71888 583986
rect 71568 583718 71610 583954
rect 71846 583718 71888 583954
rect 71568 583634 71888 583718
rect 71568 583398 71610 583634
rect 71846 583398 71888 583634
rect 71568 583366 71888 583398
rect 102288 583954 102608 583986
rect 102288 583718 102330 583954
rect 102566 583718 102608 583954
rect 102288 583634 102608 583718
rect 102288 583398 102330 583634
rect 102566 583398 102608 583634
rect 102288 583366 102608 583398
rect 133008 583954 133328 583986
rect 133008 583718 133050 583954
rect 133286 583718 133328 583954
rect 133008 583634 133328 583718
rect 133008 583398 133050 583634
rect 133286 583398 133328 583634
rect 133008 583366 133328 583398
rect 163728 583954 164048 583986
rect 163728 583718 163770 583954
rect 164006 583718 164048 583954
rect 163728 583634 164048 583718
rect 163728 583398 163770 583634
rect 164006 583398 164048 583634
rect 163728 583366 164048 583398
rect 194448 583954 194768 583986
rect 194448 583718 194490 583954
rect 194726 583718 194768 583954
rect 194448 583634 194768 583718
rect 194448 583398 194490 583634
rect 194726 583398 194768 583634
rect 194448 583366 194768 583398
rect 225168 583954 225488 583986
rect 225168 583718 225210 583954
rect 225446 583718 225488 583954
rect 225168 583634 225488 583718
rect 225168 583398 225210 583634
rect 225446 583398 225488 583634
rect 225168 583366 225488 583398
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 56208 579454 56528 579486
rect 56208 579218 56250 579454
rect 56486 579218 56528 579454
rect 56208 579134 56528 579218
rect 56208 578898 56250 579134
rect 56486 578898 56528 579134
rect 56208 578866 56528 578898
rect 86928 579454 87248 579486
rect 86928 579218 86970 579454
rect 87206 579218 87248 579454
rect 86928 579134 87248 579218
rect 86928 578898 86970 579134
rect 87206 578898 87248 579134
rect 86928 578866 87248 578898
rect 117648 579454 117968 579486
rect 117648 579218 117690 579454
rect 117926 579218 117968 579454
rect 117648 579134 117968 579218
rect 117648 578898 117690 579134
rect 117926 578898 117968 579134
rect 117648 578866 117968 578898
rect 148368 579454 148688 579486
rect 148368 579218 148410 579454
rect 148646 579218 148688 579454
rect 148368 579134 148688 579218
rect 148368 578898 148410 579134
rect 148646 578898 148688 579134
rect 148368 578866 148688 578898
rect 179088 579454 179408 579486
rect 179088 579218 179130 579454
rect 179366 579218 179408 579454
rect 179088 579134 179408 579218
rect 179088 578898 179130 579134
rect 179366 578898 179408 579134
rect 179088 578866 179408 578898
rect 209808 579454 210128 579486
rect 209808 579218 209850 579454
rect 210086 579218 210128 579454
rect 209808 579134 210128 579218
rect 209808 578898 209850 579134
rect 210086 578898 210128 579134
rect 209808 578866 210128 578898
rect 240528 579454 240848 579486
rect 240528 579218 240570 579454
rect 240806 579218 240848 579454
rect 240528 579134 240848 579218
rect 240528 578898 240570 579134
rect 240806 578898 240848 579134
rect 240528 578866 240848 578898
rect 71568 547954 71888 547986
rect 71568 547718 71610 547954
rect 71846 547718 71888 547954
rect 71568 547634 71888 547718
rect 71568 547398 71610 547634
rect 71846 547398 71888 547634
rect 71568 547366 71888 547398
rect 102288 547954 102608 547986
rect 102288 547718 102330 547954
rect 102566 547718 102608 547954
rect 102288 547634 102608 547718
rect 102288 547398 102330 547634
rect 102566 547398 102608 547634
rect 102288 547366 102608 547398
rect 133008 547954 133328 547986
rect 133008 547718 133050 547954
rect 133286 547718 133328 547954
rect 133008 547634 133328 547718
rect 133008 547398 133050 547634
rect 133286 547398 133328 547634
rect 133008 547366 133328 547398
rect 163728 547954 164048 547986
rect 163728 547718 163770 547954
rect 164006 547718 164048 547954
rect 163728 547634 164048 547718
rect 163728 547398 163770 547634
rect 164006 547398 164048 547634
rect 163728 547366 164048 547398
rect 194448 547954 194768 547986
rect 194448 547718 194490 547954
rect 194726 547718 194768 547954
rect 194448 547634 194768 547718
rect 194448 547398 194490 547634
rect 194726 547398 194768 547634
rect 194448 547366 194768 547398
rect 225168 547954 225488 547986
rect 225168 547718 225210 547954
rect 225446 547718 225488 547954
rect 225168 547634 225488 547718
rect 225168 547398 225210 547634
rect 225446 547398 225488 547634
rect 225168 547366 225488 547398
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 56208 543454 56528 543486
rect 56208 543218 56250 543454
rect 56486 543218 56528 543454
rect 56208 543134 56528 543218
rect 56208 542898 56250 543134
rect 56486 542898 56528 543134
rect 56208 542866 56528 542898
rect 86928 543454 87248 543486
rect 86928 543218 86970 543454
rect 87206 543218 87248 543454
rect 86928 543134 87248 543218
rect 86928 542898 86970 543134
rect 87206 542898 87248 543134
rect 86928 542866 87248 542898
rect 117648 543454 117968 543486
rect 117648 543218 117690 543454
rect 117926 543218 117968 543454
rect 117648 543134 117968 543218
rect 117648 542898 117690 543134
rect 117926 542898 117968 543134
rect 117648 542866 117968 542898
rect 148368 543454 148688 543486
rect 148368 543218 148410 543454
rect 148646 543218 148688 543454
rect 148368 543134 148688 543218
rect 148368 542898 148410 543134
rect 148646 542898 148688 543134
rect 148368 542866 148688 542898
rect 179088 543454 179408 543486
rect 179088 543218 179130 543454
rect 179366 543218 179408 543454
rect 179088 543134 179408 543218
rect 179088 542898 179130 543134
rect 179366 542898 179408 543134
rect 179088 542866 179408 542898
rect 209808 543454 210128 543486
rect 209808 543218 209850 543454
rect 210086 543218 210128 543454
rect 209808 543134 210128 543218
rect 209808 542898 209850 543134
rect 210086 542898 210128 543134
rect 209808 542866 210128 542898
rect 240528 543454 240848 543486
rect 240528 543218 240570 543454
rect 240806 543218 240848 543454
rect 240528 543134 240848 543218
rect 240528 542898 240570 543134
rect 240806 542898 240848 543134
rect 240528 542866 240848 542898
rect 71568 511954 71888 511986
rect 71568 511718 71610 511954
rect 71846 511718 71888 511954
rect 71568 511634 71888 511718
rect 71568 511398 71610 511634
rect 71846 511398 71888 511634
rect 71568 511366 71888 511398
rect 102288 511954 102608 511986
rect 102288 511718 102330 511954
rect 102566 511718 102608 511954
rect 102288 511634 102608 511718
rect 102288 511398 102330 511634
rect 102566 511398 102608 511634
rect 102288 511366 102608 511398
rect 133008 511954 133328 511986
rect 133008 511718 133050 511954
rect 133286 511718 133328 511954
rect 133008 511634 133328 511718
rect 133008 511398 133050 511634
rect 133286 511398 133328 511634
rect 133008 511366 133328 511398
rect 163728 511954 164048 511986
rect 163728 511718 163770 511954
rect 164006 511718 164048 511954
rect 163728 511634 164048 511718
rect 163728 511398 163770 511634
rect 164006 511398 164048 511634
rect 163728 511366 164048 511398
rect 194448 511954 194768 511986
rect 194448 511718 194490 511954
rect 194726 511718 194768 511954
rect 194448 511634 194768 511718
rect 194448 511398 194490 511634
rect 194726 511398 194768 511634
rect 194448 511366 194768 511398
rect 225168 511954 225488 511986
rect 225168 511718 225210 511954
rect 225446 511718 225488 511954
rect 225168 511634 225488 511718
rect 225168 511398 225210 511634
rect 225446 511398 225488 511634
rect 225168 511366 225488 511398
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 56208 507454 56528 507486
rect 56208 507218 56250 507454
rect 56486 507218 56528 507454
rect 56208 507134 56528 507218
rect 56208 506898 56250 507134
rect 56486 506898 56528 507134
rect 56208 506866 56528 506898
rect 86928 507454 87248 507486
rect 86928 507218 86970 507454
rect 87206 507218 87248 507454
rect 86928 507134 87248 507218
rect 86928 506898 86970 507134
rect 87206 506898 87248 507134
rect 86928 506866 87248 506898
rect 117648 507454 117968 507486
rect 117648 507218 117690 507454
rect 117926 507218 117968 507454
rect 117648 507134 117968 507218
rect 117648 506898 117690 507134
rect 117926 506898 117968 507134
rect 117648 506866 117968 506898
rect 148368 507454 148688 507486
rect 148368 507218 148410 507454
rect 148646 507218 148688 507454
rect 148368 507134 148688 507218
rect 148368 506898 148410 507134
rect 148646 506898 148688 507134
rect 148368 506866 148688 506898
rect 179088 507454 179408 507486
rect 179088 507218 179130 507454
rect 179366 507218 179408 507454
rect 179088 507134 179408 507218
rect 179088 506898 179130 507134
rect 179366 506898 179408 507134
rect 179088 506866 179408 506898
rect 209808 507454 210128 507486
rect 209808 507218 209850 507454
rect 210086 507218 210128 507454
rect 209808 507134 210128 507218
rect 209808 506898 209850 507134
rect 210086 506898 210128 507134
rect 209808 506866 210128 506898
rect 240528 507454 240848 507486
rect 240528 507218 240570 507454
rect 240806 507218 240848 507454
rect 240528 507134 240848 507218
rect 240528 506898 240570 507134
rect 240806 506898 240848 507134
rect 240528 506866 240848 506898
rect 51211 479772 51277 479773
rect 51211 479708 51212 479772
rect 51276 479708 51277 479772
rect 51211 479707 51277 479708
rect 51214 477597 51274 479707
rect 51211 477596 51277 477597
rect 51211 477532 51212 477596
rect 51276 477532 51277 477596
rect 51211 477531 51277 477532
rect 71568 475954 71888 475986
rect 71568 475718 71610 475954
rect 71846 475718 71888 475954
rect 71568 475634 71888 475718
rect 71568 475398 71610 475634
rect 71846 475398 71888 475634
rect 71568 475366 71888 475398
rect 102288 475954 102608 475986
rect 102288 475718 102330 475954
rect 102566 475718 102608 475954
rect 102288 475634 102608 475718
rect 102288 475398 102330 475634
rect 102566 475398 102608 475634
rect 102288 475366 102608 475398
rect 133008 475954 133328 475986
rect 133008 475718 133050 475954
rect 133286 475718 133328 475954
rect 133008 475634 133328 475718
rect 133008 475398 133050 475634
rect 133286 475398 133328 475634
rect 133008 475366 133328 475398
rect 163728 475954 164048 475986
rect 163728 475718 163770 475954
rect 164006 475718 164048 475954
rect 163728 475634 164048 475718
rect 163728 475398 163770 475634
rect 164006 475398 164048 475634
rect 163728 475366 164048 475398
rect 194448 475954 194768 475986
rect 194448 475718 194490 475954
rect 194726 475718 194768 475954
rect 194448 475634 194768 475718
rect 194448 475398 194490 475634
rect 194726 475398 194768 475634
rect 194448 475366 194768 475398
rect 225168 475954 225488 475986
rect 225168 475718 225210 475954
rect 225446 475718 225488 475954
rect 225168 475634 225488 475718
rect 225168 475398 225210 475634
rect 225446 475398 225488 475634
rect 225168 475366 225488 475398
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 56208 471454 56528 471486
rect 56208 471218 56250 471454
rect 56486 471218 56528 471454
rect 56208 471134 56528 471218
rect 56208 470898 56250 471134
rect 56486 470898 56528 471134
rect 56208 470866 56528 470898
rect 86928 471454 87248 471486
rect 86928 471218 86970 471454
rect 87206 471218 87248 471454
rect 86928 471134 87248 471218
rect 86928 470898 86970 471134
rect 87206 470898 87248 471134
rect 86928 470866 87248 470898
rect 117648 471454 117968 471486
rect 117648 471218 117690 471454
rect 117926 471218 117968 471454
rect 117648 471134 117968 471218
rect 117648 470898 117690 471134
rect 117926 470898 117968 471134
rect 117648 470866 117968 470898
rect 148368 471454 148688 471486
rect 148368 471218 148410 471454
rect 148646 471218 148688 471454
rect 148368 471134 148688 471218
rect 148368 470898 148410 471134
rect 148646 470898 148688 471134
rect 148368 470866 148688 470898
rect 179088 471454 179408 471486
rect 179088 471218 179130 471454
rect 179366 471218 179408 471454
rect 179088 471134 179408 471218
rect 179088 470898 179130 471134
rect 179366 470898 179408 471134
rect 179088 470866 179408 470898
rect 209808 471454 210128 471486
rect 209808 471218 209850 471454
rect 210086 471218 210128 471454
rect 209808 471134 210128 471218
rect 209808 470898 209850 471134
rect 210086 470898 210128 471134
rect 209808 470866 210128 470898
rect 240528 471454 240848 471486
rect 240528 471218 240570 471454
rect 240806 471218 240848 471454
rect 240528 471134 240848 471218
rect 240528 470898 240570 471134
rect 240806 470898 240848 471134
rect 240528 470866 240848 470898
rect 71568 439954 71888 439986
rect 71568 439718 71610 439954
rect 71846 439718 71888 439954
rect 71568 439634 71888 439718
rect 71568 439398 71610 439634
rect 71846 439398 71888 439634
rect 71568 439366 71888 439398
rect 102288 439954 102608 439986
rect 102288 439718 102330 439954
rect 102566 439718 102608 439954
rect 102288 439634 102608 439718
rect 102288 439398 102330 439634
rect 102566 439398 102608 439634
rect 102288 439366 102608 439398
rect 133008 439954 133328 439986
rect 133008 439718 133050 439954
rect 133286 439718 133328 439954
rect 133008 439634 133328 439718
rect 133008 439398 133050 439634
rect 133286 439398 133328 439634
rect 133008 439366 133328 439398
rect 163728 439954 164048 439986
rect 163728 439718 163770 439954
rect 164006 439718 164048 439954
rect 163728 439634 164048 439718
rect 163728 439398 163770 439634
rect 164006 439398 164048 439634
rect 163728 439366 164048 439398
rect 194448 439954 194768 439986
rect 194448 439718 194490 439954
rect 194726 439718 194768 439954
rect 194448 439634 194768 439718
rect 194448 439398 194490 439634
rect 194726 439398 194768 439634
rect 194448 439366 194768 439398
rect 225168 439954 225488 439986
rect 225168 439718 225210 439954
rect 225446 439718 225488 439954
rect 225168 439634 225488 439718
rect 225168 439398 225210 439634
rect 225446 439398 225488 439634
rect 225168 439366 225488 439398
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 56208 435454 56528 435486
rect 56208 435218 56250 435454
rect 56486 435218 56528 435454
rect 56208 435134 56528 435218
rect 56208 434898 56250 435134
rect 56486 434898 56528 435134
rect 56208 434866 56528 434898
rect 86928 435454 87248 435486
rect 86928 435218 86970 435454
rect 87206 435218 87248 435454
rect 86928 435134 87248 435218
rect 86928 434898 86970 435134
rect 87206 434898 87248 435134
rect 86928 434866 87248 434898
rect 117648 435454 117968 435486
rect 117648 435218 117690 435454
rect 117926 435218 117968 435454
rect 117648 435134 117968 435218
rect 117648 434898 117690 435134
rect 117926 434898 117968 435134
rect 117648 434866 117968 434898
rect 148368 435454 148688 435486
rect 148368 435218 148410 435454
rect 148646 435218 148688 435454
rect 148368 435134 148688 435218
rect 148368 434898 148410 435134
rect 148646 434898 148688 435134
rect 148368 434866 148688 434898
rect 179088 435454 179408 435486
rect 179088 435218 179130 435454
rect 179366 435218 179408 435454
rect 179088 435134 179408 435218
rect 179088 434898 179130 435134
rect 179366 434898 179408 435134
rect 179088 434866 179408 434898
rect 209808 435454 210128 435486
rect 209808 435218 209850 435454
rect 210086 435218 210128 435454
rect 209808 435134 210128 435218
rect 209808 434898 209850 435134
rect 210086 434898 210128 435134
rect 209808 434866 210128 434898
rect 240528 435454 240848 435486
rect 240528 435218 240570 435454
rect 240806 435218 240848 435454
rect 240528 435134 240848 435218
rect 240528 434898 240570 435134
rect 240806 434898 240848 435134
rect 240528 434866 240848 434898
rect 71568 403954 71888 403986
rect 71568 403718 71610 403954
rect 71846 403718 71888 403954
rect 71568 403634 71888 403718
rect 71568 403398 71610 403634
rect 71846 403398 71888 403634
rect 71568 403366 71888 403398
rect 102288 403954 102608 403986
rect 102288 403718 102330 403954
rect 102566 403718 102608 403954
rect 102288 403634 102608 403718
rect 102288 403398 102330 403634
rect 102566 403398 102608 403634
rect 102288 403366 102608 403398
rect 133008 403954 133328 403986
rect 133008 403718 133050 403954
rect 133286 403718 133328 403954
rect 133008 403634 133328 403718
rect 133008 403398 133050 403634
rect 133286 403398 133328 403634
rect 133008 403366 133328 403398
rect 163728 403954 164048 403986
rect 163728 403718 163770 403954
rect 164006 403718 164048 403954
rect 163728 403634 164048 403718
rect 163728 403398 163770 403634
rect 164006 403398 164048 403634
rect 163728 403366 164048 403398
rect 194448 403954 194768 403986
rect 194448 403718 194490 403954
rect 194726 403718 194768 403954
rect 194448 403634 194768 403718
rect 194448 403398 194490 403634
rect 194726 403398 194768 403634
rect 194448 403366 194768 403398
rect 225168 403954 225488 403986
rect 225168 403718 225210 403954
rect 225446 403718 225488 403954
rect 225168 403634 225488 403718
rect 225168 403398 225210 403634
rect 225446 403398 225488 403634
rect 225168 403366 225488 403398
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 56208 399454 56528 399486
rect 56208 399218 56250 399454
rect 56486 399218 56528 399454
rect 56208 399134 56528 399218
rect 56208 398898 56250 399134
rect 56486 398898 56528 399134
rect 56208 398866 56528 398898
rect 86928 399454 87248 399486
rect 86928 399218 86970 399454
rect 87206 399218 87248 399454
rect 86928 399134 87248 399218
rect 86928 398898 86970 399134
rect 87206 398898 87248 399134
rect 86928 398866 87248 398898
rect 117648 399454 117968 399486
rect 117648 399218 117690 399454
rect 117926 399218 117968 399454
rect 117648 399134 117968 399218
rect 117648 398898 117690 399134
rect 117926 398898 117968 399134
rect 117648 398866 117968 398898
rect 148368 399454 148688 399486
rect 148368 399218 148410 399454
rect 148646 399218 148688 399454
rect 148368 399134 148688 399218
rect 148368 398898 148410 399134
rect 148646 398898 148688 399134
rect 148368 398866 148688 398898
rect 179088 399454 179408 399486
rect 179088 399218 179130 399454
rect 179366 399218 179408 399454
rect 179088 399134 179408 399218
rect 179088 398898 179130 399134
rect 179366 398898 179408 399134
rect 179088 398866 179408 398898
rect 209808 399454 210128 399486
rect 209808 399218 209850 399454
rect 210086 399218 210128 399454
rect 209808 399134 210128 399218
rect 209808 398898 209850 399134
rect 210086 398898 210128 399134
rect 209808 398866 210128 398898
rect 240528 399454 240848 399486
rect 240528 399218 240570 399454
rect 240806 399218 240848 399454
rect 240528 399134 240848 399218
rect 240528 398898 240570 399134
rect 240806 398898 240848 399134
rect 240528 398866 240848 398898
rect 71568 367954 71888 367986
rect 71568 367718 71610 367954
rect 71846 367718 71888 367954
rect 71568 367634 71888 367718
rect 71568 367398 71610 367634
rect 71846 367398 71888 367634
rect 71568 367366 71888 367398
rect 102288 367954 102608 367986
rect 102288 367718 102330 367954
rect 102566 367718 102608 367954
rect 102288 367634 102608 367718
rect 102288 367398 102330 367634
rect 102566 367398 102608 367634
rect 102288 367366 102608 367398
rect 133008 367954 133328 367986
rect 133008 367718 133050 367954
rect 133286 367718 133328 367954
rect 133008 367634 133328 367718
rect 133008 367398 133050 367634
rect 133286 367398 133328 367634
rect 133008 367366 133328 367398
rect 163728 367954 164048 367986
rect 163728 367718 163770 367954
rect 164006 367718 164048 367954
rect 163728 367634 164048 367718
rect 163728 367398 163770 367634
rect 164006 367398 164048 367634
rect 163728 367366 164048 367398
rect 194448 367954 194768 367986
rect 194448 367718 194490 367954
rect 194726 367718 194768 367954
rect 194448 367634 194768 367718
rect 194448 367398 194490 367634
rect 194726 367398 194768 367634
rect 194448 367366 194768 367398
rect 225168 367954 225488 367986
rect 225168 367718 225210 367954
rect 225446 367718 225488 367954
rect 225168 367634 225488 367718
rect 225168 367398 225210 367634
rect 225446 367398 225488 367634
rect 225168 367366 225488 367398
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 56208 363454 56528 363486
rect 56208 363218 56250 363454
rect 56486 363218 56528 363454
rect 56208 363134 56528 363218
rect 56208 362898 56250 363134
rect 56486 362898 56528 363134
rect 56208 362866 56528 362898
rect 86928 363454 87248 363486
rect 86928 363218 86970 363454
rect 87206 363218 87248 363454
rect 86928 363134 87248 363218
rect 86928 362898 86970 363134
rect 87206 362898 87248 363134
rect 86928 362866 87248 362898
rect 117648 363454 117968 363486
rect 117648 363218 117690 363454
rect 117926 363218 117968 363454
rect 117648 363134 117968 363218
rect 117648 362898 117690 363134
rect 117926 362898 117968 363134
rect 117648 362866 117968 362898
rect 148368 363454 148688 363486
rect 148368 363218 148410 363454
rect 148646 363218 148688 363454
rect 148368 363134 148688 363218
rect 148368 362898 148410 363134
rect 148646 362898 148688 363134
rect 148368 362866 148688 362898
rect 179088 363454 179408 363486
rect 179088 363218 179130 363454
rect 179366 363218 179408 363454
rect 179088 363134 179408 363218
rect 179088 362898 179130 363134
rect 179366 362898 179408 363134
rect 179088 362866 179408 362898
rect 209808 363454 210128 363486
rect 209808 363218 209850 363454
rect 210086 363218 210128 363454
rect 209808 363134 210128 363218
rect 209808 362898 209850 363134
rect 210086 362898 210128 363134
rect 209808 362866 210128 362898
rect 240528 363454 240848 363486
rect 240528 363218 240570 363454
rect 240806 363218 240848 363454
rect 240528 363134 240848 363218
rect 240528 362898 240570 363134
rect 240806 362898 240848 363134
rect 240528 362866 240848 362898
rect 71568 331954 71888 331986
rect 71568 331718 71610 331954
rect 71846 331718 71888 331954
rect 71568 331634 71888 331718
rect 71568 331398 71610 331634
rect 71846 331398 71888 331634
rect 71568 331366 71888 331398
rect 102288 331954 102608 331986
rect 102288 331718 102330 331954
rect 102566 331718 102608 331954
rect 102288 331634 102608 331718
rect 102288 331398 102330 331634
rect 102566 331398 102608 331634
rect 102288 331366 102608 331398
rect 133008 331954 133328 331986
rect 133008 331718 133050 331954
rect 133286 331718 133328 331954
rect 133008 331634 133328 331718
rect 133008 331398 133050 331634
rect 133286 331398 133328 331634
rect 133008 331366 133328 331398
rect 163728 331954 164048 331986
rect 163728 331718 163770 331954
rect 164006 331718 164048 331954
rect 163728 331634 164048 331718
rect 163728 331398 163770 331634
rect 164006 331398 164048 331634
rect 163728 331366 164048 331398
rect 194448 331954 194768 331986
rect 194448 331718 194490 331954
rect 194726 331718 194768 331954
rect 194448 331634 194768 331718
rect 194448 331398 194490 331634
rect 194726 331398 194768 331634
rect 194448 331366 194768 331398
rect 225168 331954 225488 331986
rect 225168 331718 225210 331954
rect 225446 331718 225488 331954
rect 225168 331634 225488 331718
rect 225168 331398 225210 331634
rect 225446 331398 225488 331634
rect 225168 331366 225488 331398
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 56208 327454 56528 327486
rect 56208 327218 56250 327454
rect 56486 327218 56528 327454
rect 56208 327134 56528 327218
rect 56208 326898 56250 327134
rect 56486 326898 56528 327134
rect 56208 326866 56528 326898
rect 86928 327454 87248 327486
rect 86928 327218 86970 327454
rect 87206 327218 87248 327454
rect 86928 327134 87248 327218
rect 86928 326898 86970 327134
rect 87206 326898 87248 327134
rect 86928 326866 87248 326898
rect 117648 327454 117968 327486
rect 117648 327218 117690 327454
rect 117926 327218 117968 327454
rect 117648 327134 117968 327218
rect 117648 326898 117690 327134
rect 117926 326898 117968 327134
rect 117648 326866 117968 326898
rect 148368 327454 148688 327486
rect 148368 327218 148410 327454
rect 148646 327218 148688 327454
rect 148368 327134 148688 327218
rect 148368 326898 148410 327134
rect 148646 326898 148688 327134
rect 148368 326866 148688 326898
rect 179088 327454 179408 327486
rect 179088 327218 179130 327454
rect 179366 327218 179408 327454
rect 179088 327134 179408 327218
rect 179088 326898 179130 327134
rect 179366 326898 179408 327134
rect 179088 326866 179408 326898
rect 209808 327454 210128 327486
rect 209808 327218 209850 327454
rect 210086 327218 210128 327454
rect 209808 327134 210128 327218
rect 209808 326898 209850 327134
rect 210086 326898 210128 327134
rect 209808 326866 210128 326898
rect 240528 327454 240848 327486
rect 240528 327218 240570 327454
rect 240806 327218 240848 327454
rect 240528 327134 240848 327218
rect 240528 326898 240570 327134
rect 240806 326898 240848 327134
rect 240528 326866 240848 326898
rect 71568 295954 71888 295986
rect 71568 295718 71610 295954
rect 71846 295718 71888 295954
rect 71568 295634 71888 295718
rect 71568 295398 71610 295634
rect 71846 295398 71888 295634
rect 71568 295366 71888 295398
rect 102288 295954 102608 295986
rect 102288 295718 102330 295954
rect 102566 295718 102608 295954
rect 102288 295634 102608 295718
rect 102288 295398 102330 295634
rect 102566 295398 102608 295634
rect 102288 295366 102608 295398
rect 133008 295954 133328 295986
rect 133008 295718 133050 295954
rect 133286 295718 133328 295954
rect 133008 295634 133328 295718
rect 133008 295398 133050 295634
rect 133286 295398 133328 295634
rect 133008 295366 133328 295398
rect 163728 295954 164048 295986
rect 163728 295718 163770 295954
rect 164006 295718 164048 295954
rect 163728 295634 164048 295718
rect 163728 295398 163770 295634
rect 164006 295398 164048 295634
rect 163728 295366 164048 295398
rect 194448 295954 194768 295986
rect 194448 295718 194490 295954
rect 194726 295718 194768 295954
rect 194448 295634 194768 295718
rect 194448 295398 194490 295634
rect 194726 295398 194768 295634
rect 194448 295366 194768 295398
rect 225168 295954 225488 295986
rect 225168 295718 225210 295954
rect 225446 295718 225488 295954
rect 225168 295634 225488 295718
rect 225168 295398 225210 295634
rect 225446 295398 225488 295634
rect 225168 295366 225488 295398
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 56208 291454 56528 291486
rect 56208 291218 56250 291454
rect 56486 291218 56528 291454
rect 56208 291134 56528 291218
rect 56208 290898 56250 291134
rect 56486 290898 56528 291134
rect 56208 290866 56528 290898
rect 86928 291454 87248 291486
rect 86928 291218 86970 291454
rect 87206 291218 87248 291454
rect 86928 291134 87248 291218
rect 86928 290898 86970 291134
rect 87206 290898 87248 291134
rect 86928 290866 87248 290898
rect 117648 291454 117968 291486
rect 117648 291218 117690 291454
rect 117926 291218 117968 291454
rect 117648 291134 117968 291218
rect 117648 290898 117690 291134
rect 117926 290898 117968 291134
rect 117648 290866 117968 290898
rect 148368 291454 148688 291486
rect 148368 291218 148410 291454
rect 148646 291218 148688 291454
rect 148368 291134 148688 291218
rect 148368 290898 148410 291134
rect 148646 290898 148688 291134
rect 148368 290866 148688 290898
rect 179088 291454 179408 291486
rect 179088 291218 179130 291454
rect 179366 291218 179408 291454
rect 179088 291134 179408 291218
rect 179088 290898 179130 291134
rect 179366 290898 179408 291134
rect 179088 290866 179408 290898
rect 209808 291454 210128 291486
rect 209808 291218 209850 291454
rect 210086 291218 210128 291454
rect 209808 291134 210128 291218
rect 209808 290898 209850 291134
rect 210086 290898 210128 291134
rect 209808 290866 210128 290898
rect 240528 291454 240848 291486
rect 240528 291218 240570 291454
rect 240806 291218 240848 291454
rect 240528 291134 240848 291218
rect 240528 290898 240570 291134
rect 240806 290898 240848 291134
rect 240528 290866 240848 290898
rect 51294 268954 51914 278000
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 49555 223548 49621 223549
rect 49555 223484 49556 223548
rect 49620 223484 49621 223548
rect 49555 223483 49621 223484
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 196954 51914 232398
rect 55794 273454 56414 278000
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 222000 56414 236898
rect 60294 277954 60914 278000
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 222000 60914 241398
rect 78294 259954 78914 278000
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 222000 78914 223398
rect 82794 264454 83414 278000
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 222000 83414 227898
rect 87294 268954 87914 278000
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 222000 87914 232398
rect 91794 273454 92414 278000
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 222000 92414 236898
rect 96294 277954 96914 278000
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 222000 96914 241398
rect 114294 259954 114914 278000
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 222000 114914 223398
rect 118794 264454 119414 278000
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 222000 119414 227898
rect 123294 268954 123914 278000
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 222000 123914 232398
rect 127794 273454 128414 278000
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 222000 128414 236898
rect 132294 277954 132914 278000
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 222000 132914 241398
rect 150294 259954 150914 278000
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 222000 150914 223398
rect 154794 264454 155414 278000
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 222000 155414 227898
rect 159294 268954 159914 278000
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 222000 159914 232398
rect 163794 273454 164414 278000
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 222000 164414 236898
rect 168294 277954 168914 278000
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 222000 168914 241398
rect 186294 259954 186914 278000
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 222000 186914 223398
rect 190794 264454 191414 278000
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 222000 191414 227898
rect 195294 268954 195914 278000
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 222000 195914 232398
rect 199794 273454 200414 278000
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 222000 200414 236898
rect 204294 277954 204914 278000
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 222000 204914 241398
rect 222294 259954 222914 278000
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 222000 222914 223398
rect 226794 264454 227414 278000
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 57835 218652 57901 218653
rect 57835 218588 57836 218652
rect 57900 218588 57901 218652
rect 57835 218587 57901 218588
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 57838 131749 57898 218587
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 79568 187954 79888 187986
rect 79568 187718 79610 187954
rect 79846 187718 79888 187954
rect 79568 187634 79888 187718
rect 79568 187398 79610 187634
rect 79846 187398 79888 187634
rect 79568 187366 79888 187398
rect 110288 187954 110608 187986
rect 110288 187718 110330 187954
rect 110566 187718 110608 187954
rect 110288 187634 110608 187718
rect 110288 187398 110330 187634
rect 110566 187398 110608 187634
rect 110288 187366 110608 187398
rect 141008 187954 141328 187986
rect 141008 187718 141050 187954
rect 141286 187718 141328 187954
rect 141008 187634 141328 187718
rect 141008 187398 141050 187634
rect 141286 187398 141328 187634
rect 141008 187366 141328 187398
rect 171728 187954 172048 187986
rect 171728 187718 171770 187954
rect 172006 187718 172048 187954
rect 171728 187634 172048 187718
rect 171728 187398 171770 187634
rect 172006 187398 172048 187634
rect 171728 187366 172048 187398
rect 202448 187954 202768 187986
rect 202448 187718 202490 187954
rect 202726 187718 202768 187954
rect 202448 187634 202768 187718
rect 202448 187398 202490 187634
rect 202726 187398 202768 187634
rect 202448 187366 202768 187398
rect 64208 183454 64528 183486
rect 64208 183218 64250 183454
rect 64486 183218 64528 183454
rect 64208 183134 64528 183218
rect 64208 182898 64250 183134
rect 64486 182898 64528 183134
rect 64208 182866 64528 182898
rect 94928 183454 95248 183486
rect 94928 183218 94970 183454
rect 95206 183218 95248 183454
rect 94928 183134 95248 183218
rect 94928 182898 94970 183134
rect 95206 182898 95248 183134
rect 94928 182866 95248 182898
rect 125648 183454 125968 183486
rect 125648 183218 125690 183454
rect 125926 183218 125968 183454
rect 125648 183134 125968 183218
rect 125648 182898 125690 183134
rect 125926 182898 125968 183134
rect 125648 182866 125968 182898
rect 156368 183454 156688 183486
rect 156368 183218 156410 183454
rect 156646 183218 156688 183454
rect 156368 183134 156688 183218
rect 156368 182898 156410 183134
rect 156646 182898 156688 183134
rect 156368 182866 156688 182898
rect 187088 183454 187408 183486
rect 187088 183218 187130 183454
rect 187366 183218 187408 183454
rect 187088 183134 187408 183218
rect 187088 182898 187130 183134
rect 187366 182898 187408 183134
rect 187088 182866 187408 182898
rect 217808 183454 218128 183486
rect 217808 183218 217850 183454
rect 218086 183218 218128 183454
rect 217808 183134 218128 183218
rect 217808 182898 217850 183134
rect 218086 182898 218128 183134
rect 217808 182866 218128 182898
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 79568 151954 79888 151986
rect 79568 151718 79610 151954
rect 79846 151718 79888 151954
rect 79568 151634 79888 151718
rect 79568 151398 79610 151634
rect 79846 151398 79888 151634
rect 79568 151366 79888 151398
rect 110288 151954 110608 151986
rect 110288 151718 110330 151954
rect 110566 151718 110608 151954
rect 110288 151634 110608 151718
rect 110288 151398 110330 151634
rect 110566 151398 110608 151634
rect 110288 151366 110608 151398
rect 141008 151954 141328 151986
rect 141008 151718 141050 151954
rect 141286 151718 141328 151954
rect 141008 151634 141328 151718
rect 141008 151398 141050 151634
rect 141286 151398 141328 151634
rect 141008 151366 141328 151398
rect 171728 151954 172048 151986
rect 171728 151718 171770 151954
rect 172006 151718 172048 151954
rect 171728 151634 172048 151718
rect 171728 151398 171770 151634
rect 172006 151398 172048 151634
rect 171728 151366 172048 151398
rect 202448 151954 202768 151986
rect 202448 151718 202490 151954
rect 202726 151718 202768 151954
rect 202448 151634 202768 151718
rect 202448 151398 202490 151634
rect 202726 151398 202768 151634
rect 202448 151366 202768 151398
rect 64208 147454 64528 147486
rect 64208 147218 64250 147454
rect 64486 147218 64528 147454
rect 64208 147134 64528 147218
rect 64208 146898 64250 147134
rect 64486 146898 64528 147134
rect 64208 146866 64528 146898
rect 94928 147454 95248 147486
rect 94928 147218 94970 147454
rect 95206 147218 95248 147454
rect 94928 147134 95248 147218
rect 94928 146898 94970 147134
rect 95206 146898 95248 147134
rect 94928 146866 95248 146898
rect 125648 147454 125968 147486
rect 125648 147218 125690 147454
rect 125926 147218 125968 147454
rect 125648 147134 125968 147218
rect 125648 146898 125690 147134
rect 125926 146898 125968 147134
rect 125648 146866 125968 146898
rect 156368 147454 156688 147486
rect 156368 147218 156410 147454
rect 156646 147218 156688 147454
rect 156368 147134 156688 147218
rect 156368 146898 156410 147134
rect 156646 146898 156688 147134
rect 156368 146866 156688 146898
rect 187088 147454 187408 147486
rect 187088 147218 187130 147454
rect 187366 147218 187408 147454
rect 187088 147134 187408 147218
rect 187088 146898 187130 147134
rect 187366 146898 187408 147134
rect 187088 146866 187408 146898
rect 217808 147454 218128 147486
rect 217808 147218 217850 147454
rect 218086 147218 218128 147454
rect 217808 147134 218128 147218
rect 217808 146898 217850 147134
rect 218086 146898 218128 147134
rect 217808 146866 218128 146898
rect 57835 131748 57901 131749
rect 57835 131684 57836 131748
rect 57900 131684 57901 131748
rect 57835 131683 57901 131684
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 79568 115954 79888 115986
rect 79568 115718 79610 115954
rect 79846 115718 79888 115954
rect 79568 115634 79888 115718
rect 79568 115398 79610 115634
rect 79846 115398 79888 115634
rect 79568 115366 79888 115398
rect 110288 115954 110608 115986
rect 110288 115718 110330 115954
rect 110566 115718 110608 115954
rect 110288 115634 110608 115718
rect 110288 115398 110330 115634
rect 110566 115398 110608 115634
rect 110288 115366 110608 115398
rect 141008 115954 141328 115986
rect 141008 115718 141050 115954
rect 141286 115718 141328 115954
rect 141008 115634 141328 115718
rect 141008 115398 141050 115634
rect 141286 115398 141328 115634
rect 141008 115366 141328 115398
rect 171728 115954 172048 115986
rect 171728 115718 171770 115954
rect 172006 115718 172048 115954
rect 171728 115634 172048 115718
rect 171728 115398 171770 115634
rect 172006 115398 172048 115634
rect 171728 115366 172048 115398
rect 202448 115954 202768 115986
rect 202448 115718 202490 115954
rect 202726 115718 202768 115954
rect 202448 115634 202768 115718
rect 202448 115398 202490 115634
rect 202726 115398 202768 115634
rect 202448 115366 202768 115398
rect 64208 111454 64528 111486
rect 64208 111218 64250 111454
rect 64486 111218 64528 111454
rect 64208 111134 64528 111218
rect 64208 110898 64250 111134
rect 64486 110898 64528 111134
rect 64208 110866 64528 110898
rect 94928 111454 95248 111486
rect 94928 111218 94970 111454
rect 95206 111218 95248 111454
rect 94928 111134 95248 111218
rect 94928 110898 94970 111134
rect 95206 110898 95248 111134
rect 94928 110866 95248 110898
rect 125648 111454 125968 111486
rect 125648 111218 125690 111454
rect 125926 111218 125968 111454
rect 125648 111134 125968 111218
rect 125648 110898 125690 111134
rect 125926 110898 125968 111134
rect 125648 110866 125968 110898
rect 156368 111454 156688 111486
rect 156368 111218 156410 111454
rect 156646 111218 156688 111454
rect 156368 111134 156688 111218
rect 156368 110898 156410 111134
rect 156646 110898 156688 111134
rect 156368 110866 156688 110898
rect 187088 111454 187408 111486
rect 187088 111218 187130 111454
rect 187366 111218 187408 111454
rect 187088 111134 187408 111218
rect 187088 110898 187130 111134
rect 187366 110898 187408 111134
rect 187088 110866 187408 110898
rect 217808 111454 218128 111486
rect 217808 111218 217850 111454
rect 218086 111218 218128 111454
rect 217808 111134 218128 111218
rect 217808 110898 217850 111134
rect 218086 110898 218128 111134
rect 217808 110866 218128 110898
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 79568 79954 79888 79986
rect 79568 79718 79610 79954
rect 79846 79718 79888 79954
rect 79568 79634 79888 79718
rect 79568 79398 79610 79634
rect 79846 79398 79888 79634
rect 79568 79366 79888 79398
rect 110288 79954 110608 79986
rect 110288 79718 110330 79954
rect 110566 79718 110608 79954
rect 110288 79634 110608 79718
rect 110288 79398 110330 79634
rect 110566 79398 110608 79634
rect 110288 79366 110608 79398
rect 141008 79954 141328 79986
rect 141008 79718 141050 79954
rect 141286 79718 141328 79954
rect 141008 79634 141328 79718
rect 141008 79398 141050 79634
rect 141286 79398 141328 79634
rect 141008 79366 141328 79398
rect 171728 79954 172048 79986
rect 171728 79718 171770 79954
rect 172006 79718 172048 79954
rect 171728 79634 172048 79718
rect 171728 79398 171770 79634
rect 172006 79398 172048 79634
rect 171728 79366 172048 79398
rect 202448 79954 202768 79986
rect 202448 79718 202490 79954
rect 202726 79718 202768 79954
rect 202448 79634 202768 79718
rect 202448 79398 202490 79634
rect 202726 79398 202768 79634
rect 202448 79366 202768 79398
rect 64208 75454 64528 75486
rect 64208 75218 64250 75454
rect 64486 75218 64528 75454
rect 64208 75134 64528 75218
rect 64208 74898 64250 75134
rect 64486 74898 64528 75134
rect 64208 74866 64528 74898
rect 94928 75454 95248 75486
rect 94928 75218 94970 75454
rect 95206 75218 95248 75454
rect 94928 75134 95248 75218
rect 94928 74898 94970 75134
rect 95206 74898 95248 75134
rect 94928 74866 95248 74898
rect 125648 75454 125968 75486
rect 125648 75218 125690 75454
rect 125926 75218 125968 75454
rect 125648 75134 125968 75218
rect 125648 74898 125690 75134
rect 125926 74898 125968 75134
rect 125648 74866 125968 74898
rect 156368 75454 156688 75486
rect 156368 75218 156410 75454
rect 156646 75218 156688 75454
rect 156368 75134 156688 75218
rect 156368 74898 156410 75134
rect 156646 74898 156688 75134
rect 156368 74866 156688 74898
rect 187088 75454 187408 75486
rect 187088 75218 187130 75454
rect 187366 75218 187408 75454
rect 187088 75134 187408 75218
rect 187088 74898 187130 75134
rect 187366 74898 187408 75134
rect 187088 74866 187408 74898
rect 217808 75454 218128 75486
rect 217808 75218 217850 75454
rect 218086 75218 218128 75454
rect 217808 75134 218128 75218
rect 217808 74898 217850 75134
rect 218086 74898 218128 75134
rect 217808 74866 218128 74898
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 57454 56414 58000
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 25954 60914 58000
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 30454 65414 58000
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 34954 69914 58000
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 43954 78914 58000
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 48454 83414 58000
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 52954 87914 58000
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 25954 96914 58000
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 30454 101414 58000
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 34954 105914 58000
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 58000
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 58000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 58000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 25954 132914 58000
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 30454 137414 58000
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 34954 141914 58000
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 43954 150914 58000
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 48454 155414 58000
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 52954 159914 58000
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 25954 168914 58000
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 30454 173414 58000
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 34954 177914 58000
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 58000
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 58000
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 52954 195914 58000
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 25954 204914 58000
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 30454 209414 58000
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 34954 213914 58000
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 43954 222914 58000
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 268954 231914 278000
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 273454 236414 278000
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 277954 240914 278000
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 246454 245414 278000
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 250954 249914 278000
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 255454 254414 278000
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 642000 276914 673398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 279371 670716 279437 670717
rect 279371 670652 279372 670716
rect 279436 670652 279437 670716
rect 279371 670651 279437 670652
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 279374 567901 279434 670651
rect 280794 642361 281414 677898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 283419 663236 283485 663237
rect 283419 663172 283420 663236
rect 283484 663172 283485 663236
rect 283419 663171 283485 663172
rect 280794 642125 280826 642361
rect 281062 642125 281146 642361
rect 281382 642125 281414 642361
rect 280794 642000 281414 642125
rect 282683 639300 282749 639301
rect 282683 639236 282684 639300
rect 282748 639236 282749 639300
rect 282683 639235 282749 639236
rect 282686 579053 282746 639235
rect 282683 579052 282749 579053
rect 282683 578988 282684 579052
rect 282748 578988 282749 579052
rect 282683 578987 282749 578988
rect 279371 567900 279437 567901
rect 279371 567836 279372 567900
rect 279436 567836 279437 567900
rect 279371 567835 279437 567836
rect 279371 564636 279437 564637
rect 279371 564572 279372 564636
rect 279436 564572 279437 564636
rect 279371 564571 279437 564572
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 493954 276914 498000
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 279374 71093 279434 564571
rect 283422 543013 283482 663171
rect 285294 646954 285914 682398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 286179 663100 286245 663101
rect 286179 663036 286180 663100
rect 286244 663036 286245 663100
rect 286179 663035 286245 663036
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 642000 285914 646398
rect 285443 639300 285509 639301
rect 285443 639236 285444 639300
rect 285508 639236 285509 639300
rect 285443 639235 285509 639236
rect 284208 615454 284528 615486
rect 284208 615218 284250 615454
rect 284486 615218 284528 615454
rect 284208 615134 284528 615218
rect 284208 614898 284250 615134
rect 284486 614898 284528 615134
rect 284208 614866 284528 614898
rect 285446 563685 285506 639235
rect 285443 563684 285509 563685
rect 285443 563620 285444 563684
rect 285508 563620 285509 563684
rect 285443 563619 285509 563620
rect 286182 543149 286242 663035
rect 289794 651454 290414 686898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 290963 661876 291029 661877
rect 290963 661812 290964 661876
rect 291028 661812 291029 661876
rect 290963 661811 291029 661812
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 642000 290414 650898
rect 288203 639300 288269 639301
rect 288203 639236 288204 639300
rect 288268 639236 288269 639300
rect 288203 639235 288269 639236
rect 289491 639300 289557 639301
rect 289491 639236 289492 639300
rect 289556 639236 289557 639300
rect 289491 639235 289557 639236
rect 288206 551445 288266 639235
rect 289494 554165 289554 639235
rect 289794 579454 290414 598000
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289491 554164 289557 554165
rect 289491 554100 289492 554164
rect 289556 554100 289557 554164
rect 289491 554099 289557 554100
rect 288203 551444 288269 551445
rect 288203 551380 288204 551444
rect 288268 551380 288269 551444
rect 288203 551379 288269 551380
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 290966 543421 291026 661811
rect 291699 660652 291765 660653
rect 291699 660588 291700 660652
rect 291764 660588 291765 660652
rect 291699 660587 291765 660588
rect 290963 543420 291029 543421
rect 290963 543356 290964 543420
rect 291028 543356 291029 543420
rect 290963 543355 291029 543356
rect 286179 543148 286245 543149
rect 286179 543084 286180 543148
rect 286244 543084 286245 543148
rect 286179 543083 286245 543084
rect 289794 543134 290414 543218
rect 283419 543012 283485 543013
rect 283419 542948 283420 543012
rect 283484 542948 283485 543012
rect 283419 542947 283485 542948
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 542000 290414 542898
rect 291702 542877 291762 660587
rect 294294 655954 294914 691398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 295931 661740 295997 661741
rect 295931 661676 295932 661740
rect 295996 661676 295997 661740
rect 295931 661675 295997 661676
rect 295011 660516 295077 660517
rect 295011 660452 295012 660516
rect 295076 660452 295077 660516
rect 295011 660451 295077 660452
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 642000 294914 655398
rect 293171 641884 293237 641885
rect 293171 641820 293172 641884
rect 293236 641820 293237 641884
rect 293171 641819 293237 641820
rect 293174 551581 293234 641819
rect 294294 583954 294914 598000
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 293171 551580 293237 551581
rect 293171 551516 293172 551580
rect 293236 551516 293237 551580
rect 293171 551515 293237 551516
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 291699 542876 291765 542877
rect 291699 542812 291700 542876
rect 291764 542812 291765 542876
rect 291699 542811 291765 542812
rect 294294 542000 294914 547398
rect 295014 542605 295074 660451
rect 295934 543285 295994 661675
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 299979 660380 300045 660381
rect 299979 660316 299980 660380
rect 300044 660316 300045 660380
rect 299979 660315 300045 660316
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 297219 659836 297285 659837
rect 297219 659772 297220 659836
rect 297284 659772 297285 659836
rect 297219 659771 297285 659772
rect 295931 543284 295997 543285
rect 295931 543220 295932 543284
rect 295996 543220 295997 543284
rect 295931 543219 295997 543220
rect 295011 542604 295077 542605
rect 295011 542540 295012 542604
rect 295076 542540 295077 542604
rect 295011 542539 295077 542540
rect 297222 542469 297282 659771
rect 298794 642000 299414 659898
rect 298323 639436 298389 639437
rect 298323 639372 298324 639436
rect 298388 639372 298389 639436
rect 298323 639371 298389 639372
rect 298326 562325 298386 639371
rect 298507 639300 298573 639301
rect 298507 639236 298508 639300
rect 298572 639236 298573 639300
rect 298507 639235 298573 639236
rect 298323 562324 298389 562325
rect 298323 562260 298324 562324
rect 298388 562260 298389 562324
rect 298323 562259 298389 562260
rect 298510 559605 298570 639235
rect 299568 619954 299888 619986
rect 299568 619718 299610 619954
rect 299846 619718 299888 619954
rect 299568 619634 299888 619718
rect 299568 619398 299610 619634
rect 299846 619398 299888 619634
rect 299568 619366 299888 619398
rect 298794 588454 299414 598000
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298507 559604 298573 559605
rect 298507 559540 298508 559604
rect 298572 559540 298573 559604
rect 298507 559539 298573 559540
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 297219 542468 297285 542469
rect 297219 542404 297220 542468
rect 297284 542404 297285 542468
rect 297219 542403 297285 542404
rect 298794 542000 299414 551898
rect 299982 542469 300042 660315
rect 303294 642000 303914 664398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 304211 661604 304277 661605
rect 304211 661540 304212 661604
rect 304276 661540 304277 661604
rect 304211 661539 304277 661540
rect 303475 639572 303541 639573
rect 303475 639508 303476 639572
rect 303540 639508 303541 639572
rect 303475 639507 303541 639508
rect 302003 639028 302069 639029
rect 302003 638964 302004 639028
rect 302068 638964 302069 639028
rect 302003 638963 302069 638964
rect 302006 600677 302066 638963
rect 303478 600677 303538 639507
rect 302003 600676 302069 600677
rect 302003 600612 302004 600676
rect 302068 600612 302069 600676
rect 302003 600611 302069 600612
rect 303475 600676 303541 600677
rect 303475 600612 303476 600676
rect 303540 600612 303541 600676
rect 303475 600611 303541 600612
rect 299979 542468 300045 542469
rect 299979 542404 299980 542468
rect 300044 542404 300045 542468
rect 299979 542403 300045 542404
rect 287283 539748 287349 539749
rect 287283 539684 287284 539748
rect 287348 539684 287349 539748
rect 287283 539683 287349 539684
rect 284891 539612 284957 539613
rect 284891 539548 284892 539612
rect 284956 539548 284957 539612
rect 284891 539547 284957 539548
rect 285995 539612 286061 539613
rect 285995 539548 285996 539612
rect 286060 539548 286061 539612
rect 285995 539547 286061 539548
rect 284208 507454 284528 507486
rect 284208 507218 284250 507454
rect 284486 507218 284528 507454
rect 284208 507134 284528 507218
rect 284208 506898 284250 507134
rect 284486 506898 284528 507134
rect 284208 506866 284528 506898
rect 280794 462454 281414 498000
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 284894 292637 284954 539547
rect 285294 466954 285914 498000
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 284891 292636 284957 292637
rect 284891 292572 284892 292636
rect 284956 292572 284957 292636
rect 284891 292571 284957 292572
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 279371 71092 279437 71093
rect 279371 71028 279372 71092
rect 279436 71028 279437 71092
rect 279371 71027 279437 71028
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285998 281893 286058 539547
rect 285995 281892 286061 281893
rect 285995 281828 285996 281892
rect 286060 281828 286061 281892
rect 285995 281827 286061 281828
rect 287286 281077 287346 539683
rect 287467 539612 287533 539613
rect 287467 539548 287468 539612
rect 287532 539548 287533 539612
rect 287467 539547 287533 539548
rect 288387 539612 288453 539613
rect 288387 539548 288388 539612
rect 288452 539548 288453 539612
rect 288387 539547 288453 539548
rect 288755 539612 288821 539613
rect 288755 539548 288756 539612
rect 288820 539548 288821 539612
rect 288755 539547 288821 539548
rect 290595 539612 290661 539613
rect 290595 539548 290596 539612
rect 290660 539548 290661 539612
rect 290595 539547 290661 539548
rect 290779 539612 290845 539613
rect 290779 539548 290780 539612
rect 290844 539548 290845 539612
rect 290779 539547 290845 539548
rect 291147 539612 291213 539613
rect 291147 539548 291148 539612
rect 291212 539548 291213 539612
rect 291147 539547 291213 539548
rect 292803 539612 292869 539613
rect 292803 539548 292804 539612
rect 292868 539548 292869 539612
rect 292803 539547 292869 539548
rect 287283 281076 287349 281077
rect 287283 281012 287284 281076
rect 287348 281012 287349 281076
rect 287283 281011 287349 281012
rect 287470 280941 287530 539547
rect 287467 280940 287533 280941
rect 287467 280876 287468 280940
rect 287532 280876 287533 280940
rect 287467 280875 287533 280876
rect 288390 280669 288450 539547
rect 288758 280805 288818 539547
rect 289794 471454 290414 498000
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 288755 280804 288821 280805
rect 288755 280740 288756 280804
rect 288820 280740 288821 280804
rect 288755 280739 288821 280740
rect 288387 280668 288453 280669
rect 288387 280604 288388 280668
rect 288452 280604 288453 280668
rect 288387 280603 288453 280604
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 255454 290414 290898
rect 290598 281213 290658 539547
rect 290782 281349 290842 539547
rect 291150 282029 291210 539547
rect 291147 282028 291213 282029
rect 291147 281964 291148 282028
rect 291212 281964 291213 282028
rect 291147 281963 291213 281964
rect 290779 281348 290845 281349
rect 290779 281284 290780 281348
rect 290844 281284 290845 281348
rect 290779 281283 290845 281284
rect 290595 281212 290661 281213
rect 290595 281148 290596 281212
rect 290660 281148 290661 281212
rect 290595 281147 290661 281148
rect 292806 280533 292866 539547
rect 299568 511954 299888 511986
rect 299568 511718 299610 511954
rect 299846 511718 299888 511954
rect 299568 511634 299888 511718
rect 299568 511398 299610 511634
rect 299846 511398 299888 511634
rect 299568 511366 299888 511398
rect 302006 499221 302066 600611
rect 303294 592954 303914 598000
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 542000 303914 556398
rect 304214 542469 304274 661539
rect 305499 661468 305565 661469
rect 305499 661404 305500 661468
rect 305564 661404 305565 661468
rect 305499 661403 305565 661404
rect 305502 542605 305562 661403
rect 307794 642000 308414 668898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 308627 661332 308693 661333
rect 308627 661268 308628 661332
rect 308692 661268 308693 661332
rect 308627 661267 308693 661268
rect 307523 640932 307589 640933
rect 307523 640868 307524 640932
rect 307588 640868 307589 640932
rect 307523 640867 307589 640868
rect 307526 600677 307586 640867
rect 307523 600676 307589 600677
rect 307523 600612 307524 600676
rect 307588 600612 307589 600676
rect 307523 600611 307589 600612
rect 307794 597454 308414 598000
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 305499 542604 305565 542605
rect 305499 542540 305500 542604
rect 305564 542540 305565 542604
rect 305499 542539 305565 542540
rect 304211 542468 304277 542469
rect 304211 542404 304212 542468
rect 304276 542404 304277 542468
rect 304211 542403 304277 542404
rect 307794 542000 308414 560898
rect 308630 542741 308690 661267
rect 309363 661196 309429 661197
rect 309363 661132 309364 661196
rect 309428 661132 309429 661196
rect 309363 661131 309429 661132
rect 309179 661060 309245 661061
rect 309179 660996 309180 661060
rect 309244 660996 309245 661060
rect 309179 660995 309245 660996
rect 308811 660244 308877 660245
rect 308811 660180 308812 660244
rect 308876 660180 308877 660244
rect 308811 660179 308877 660180
rect 308627 542740 308693 542741
rect 308627 542676 308628 542740
rect 308692 542676 308693 542740
rect 308627 542675 308693 542676
rect 308814 542469 308874 660179
rect 309182 542469 309242 660995
rect 309366 542605 309426 661131
rect 310467 660108 310533 660109
rect 310467 660044 310468 660108
rect 310532 660044 310533 660108
rect 310467 660043 310533 660044
rect 309363 542604 309429 542605
rect 309363 542540 309364 542604
rect 309428 542540 309429 542604
rect 309363 542539 309429 542540
rect 310470 542469 310530 660043
rect 311939 659972 312005 659973
rect 311939 659908 311940 659972
rect 312004 659908 312005 659972
rect 311939 659907 312005 659908
rect 311019 641748 311085 641749
rect 311019 641684 311020 641748
rect 311084 641684 311085 641748
rect 311019 641683 311085 641684
rect 311022 578917 311082 641683
rect 311019 578916 311085 578917
rect 311019 578852 311020 578916
rect 311084 578852 311085 578916
rect 311019 578851 311085 578852
rect 311942 542877 312002 659907
rect 312294 642000 312914 673398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642361 317414 677898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 317643 662964 317709 662965
rect 317643 662900 317644 662964
rect 317708 662900 317709 662964
rect 317643 662899 317709 662900
rect 316794 642125 316826 642361
rect 317062 642125 317146 642361
rect 317382 642125 317414 642361
rect 316794 642000 317414 642125
rect 314928 615454 315248 615486
rect 314928 615218 314970 615454
rect 315206 615218 315248 615454
rect 314928 615134 315248 615218
rect 314928 614898 314970 615134
rect 315206 614898 315248 615134
rect 314928 614866 315248 614898
rect 317646 543693 317706 662899
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 642000 321914 646398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 317643 543692 317709 543693
rect 317643 543628 317644 543692
rect 317708 543628 317709 543692
rect 317643 543627 317709 543628
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 311939 542876 312005 542877
rect 311939 542812 311940 542876
rect 312004 542812 312005 542876
rect 311939 542811 312005 542812
rect 308811 542468 308877 542469
rect 308811 542404 308812 542468
rect 308876 542404 308877 542468
rect 308811 542403 308877 542404
rect 309179 542468 309245 542469
rect 309179 542404 309180 542468
rect 309244 542404 309245 542468
rect 309179 542403 309245 542404
rect 310467 542468 310533 542469
rect 310467 542404 310468 542468
rect 310532 542404 310533 542468
rect 310467 542403 310533 542404
rect 314928 507454 315248 507486
rect 314928 507218 314970 507454
rect 315206 507218 315248 507454
rect 314928 507134 315248 507218
rect 314928 506898 314970 507134
rect 315206 506898 315248 507134
rect 314928 506866 315248 506898
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 302003 499220 302069 499221
rect 302003 499156 302004 499220
rect 302068 499156 302069 499220
rect 302003 499155 302069 499156
rect 294294 475954 294914 498000
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 298794 480454 299414 498000
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 303294 484954 303914 498000
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 299979 340100 300045 340101
rect 299979 340036 299980 340100
rect 300044 340036 300045 340100
rect 299979 340035 300045 340036
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298507 334660 298573 334661
rect 298507 334596 298508 334660
rect 298572 334596 298573 334660
rect 298507 334595 298573 334596
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 295931 331940 295997 331941
rect 295931 331876 295932 331940
rect 295996 331876 295997 331940
rect 295931 331875 295997 331876
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 292803 280532 292869 280533
rect 292803 280468 292804 280532
rect 292868 280468 292869 280532
rect 292803 280467 292869 280468
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 259954 294914 295398
rect 295934 282165 295994 331875
rect 297219 310044 297285 310045
rect 297219 309980 297220 310044
rect 297284 309980 297285 310044
rect 297219 309979 297285 309980
rect 295931 282164 295997 282165
rect 295931 282100 295932 282164
rect 295996 282100 295997 282164
rect 295931 282099 295997 282100
rect 297222 278085 297282 309979
rect 297219 278084 297285 278085
rect 297219 278020 297220 278084
rect 297284 278020 297285 278084
rect 297219 278019 297285 278020
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 298510 3637 298570 334595
rect 298794 332000 299414 335898
rect 299243 311404 299309 311405
rect 299243 311340 299244 311404
rect 299308 311340 299309 311404
rect 299243 311339 299309 311340
rect 299246 281485 299306 311339
rect 299243 281484 299309 281485
rect 299243 281420 299244 281484
rect 299308 281420 299309 281484
rect 299243 281419 299309 281420
rect 298794 264454 299414 278000
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 222000 299414 227898
rect 298794 48454 299414 58000
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298507 3636 298573 3637
rect 298507 3572 298508 3636
rect 298572 3572 298573 3636
rect 298507 3571 298573 3572
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 -2266 299414 11898
rect 299982 3637 300042 340035
rect 303294 332000 303914 340398
rect 307794 489454 308414 498000
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 332000 308414 344898
rect 312294 493954 312914 498000
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 332000 312914 349398
rect 316794 462454 317414 498000
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 332000 317414 353898
rect 321294 466954 321914 498000
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 332000 321914 358398
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 332000 326414 362898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 332000 330914 367398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 332000 335414 335898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 332000 339914 340398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 332000 344414 344898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 642000 357914 646398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 359411 642156 359477 642157
rect 359411 642092 359412 642156
rect 359476 642092 359477 642156
rect 359411 642091 359477 642092
rect 352794 606454 353414 641898
rect 355363 640524 355429 640525
rect 355363 640460 355364 640524
rect 355428 640460 355429 640524
rect 355363 640459 355429 640460
rect 355179 640388 355245 640389
rect 355179 640324 355180 640388
rect 355244 640324 355245 640388
rect 355179 640323 355245 640324
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 349107 518940 349173 518941
rect 349107 518876 349108 518940
rect 349172 518876 349173 518940
rect 349107 518875 349173 518876
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 332000 348914 349398
rect 300163 331260 300229 331261
rect 300163 331196 300164 331260
rect 300228 331196 300229 331260
rect 300163 331195 300229 331196
rect 300166 218245 300226 331195
rect 304208 327239 304528 327376
rect 304208 327003 304250 327239
rect 304486 327003 304528 327239
rect 304208 326866 304528 327003
rect 334928 327239 335248 327376
rect 334928 327003 334970 327239
rect 335206 327003 335248 327239
rect 334928 326866 335248 327003
rect 319568 295954 319888 295986
rect 319568 295718 319610 295954
rect 319846 295718 319888 295954
rect 319568 295634 319888 295718
rect 319568 295398 319610 295634
rect 319846 295398 319888 295634
rect 319568 295366 319888 295398
rect 304208 291454 304528 291486
rect 304208 291218 304250 291454
rect 304486 291218 304528 291454
rect 304208 291134 304528 291218
rect 304208 290898 304250 291134
rect 304486 290898 304528 291134
rect 304208 290866 304528 290898
rect 334928 291454 335248 291486
rect 334928 291218 334970 291454
rect 335206 291218 335248 291454
rect 334928 291134 335248 291218
rect 334928 290898 334970 291134
rect 335206 290898 335248 291134
rect 334928 290866 335248 290898
rect 303294 268954 303914 278000
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 222000 303914 232398
rect 307794 273454 308414 278000
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 222000 308414 236898
rect 312294 277954 312914 278000
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 222000 312914 241398
rect 330294 259954 330914 278000
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 222000 330914 223398
rect 334794 264454 335414 278000
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 222000 335414 227898
rect 339294 268954 339914 278000
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 222000 339914 232398
rect 343794 273454 344414 278000
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 222000 344414 236898
rect 348294 277954 348914 278000
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 300163 218244 300229 218245
rect 300163 218180 300164 218244
rect 300228 218180 300229 218244
rect 300163 218179 300229 218180
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 319568 187954 319888 187986
rect 319568 187718 319610 187954
rect 319846 187718 319888 187954
rect 319568 187634 319888 187718
rect 319568 187398 319610 187634
rect 319846 187398 319888 187634
rect 319568 187366 319888 187398
rect 304208 183454 304528 183486
rect 304208 183218 304250 183454
rect 304486 183218 304528 183454
rect 304208 183134 304528 183218
rect 304208 182898 304250 183134
rect 304486 182898 304528 183134
rect 304208 182866 304528 182898
rect 334928 183454 335248 183486
rect 334928 183218 334970 183454
rect 335206 183218 335248 183454
rect 334928 183134 335248 183218
rect 334928 182898 334970 183134
rect 335206 182898 335248 183134
rect 334928 182866 335248 182898
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 319568 151954 319888 151986
rect 319568 151718 319610 151954
rect 319846 151718 319888 151954
rect 319568 151634 319888 151718
rect 319568 151398 319610 151634
rect 319846 151398 319888 151634
rect 319568 151366 319888 151398
rect 304208 147454 304528 147486
rect 304208 147218 304250 147454
rect 304486 147218 304528 147454
rect 304208 147134 304528 147218
rect 304208 146898 304250 147134
rect 304486 146898 304528 147134
rect 304208 146866 304528 146898
rect 334928 147454 335248 147486
rect 334928 147218 334970 147454
rect 335206 147218 335248 147454
rect 334928 147134 335248 147218
rect 334928 146898 334970 147134
rect 335206 146898 335248 147134
rect 334928 146866 335248 146898
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 319568 115954 319888 115986
rect 319568 115718 319610 115954
rect 319846 115718 319888 115954
rect 319568 115634 319888 115718
rect 319568 115398 319610 115634
rect 319846 115398 319888 115634
rect 319568 115366 319888 115398
rect 304208 111454 304528 111486
rect 304208 111218 304250 111454
rect 304486 111218 304528 111454
rect 304208 111134 304528 111218
rect 304208 110898 304250 111134
rect 304486 110898 304528 111134
rect 304208 110866 304528 110898
rect 334928 111454 335248 111486
rect 334928 111218 334970 111454
rect 335206 111218 335248 111454
rect 334928 111134 335248 111218
rect 334928 110898 334970 111134
rect 335206 110898 335248 111134
rect 334928 110866 335248 110898
rect 340827 108356 340893 108357
rect 340827 108292 340828 108356
rect 340892 108292 340893 108356
rect 340827 108291 340893 108292
rect 340091 85508 340157 85509
rect 340091 85444 340092 85508
rect 340156 85444 340157 85508
rect 340091 85443 340157 85444
rect 319568 79954 319888 79986
rect 319568 79718 319610 79954
rect 319846 79718 319888 79954
rect 319568 79634 319888 79718
rect 319568 79398 319610 79634
rect 319846 79398 319888 79634
rect 319568 79366 319888 79398
rect 304208 75454 304528 75486
rect 304208 75218 304250 75454
rect 304486 75218 304528 75454
rect 304208 75134 304528 75218
rect 304208 74898 304250 75134
rect 304486 74898 304528 75134
rect 304208 74866 304528 74898
rect 334928 75454 335248 75486
rect 334928 75218 334970 75454
rect 335206 75218 335248 75454
rect 334928 75134 335248 75218
rect 334928 74898 334970 75134
rect 335206 74898 335248 75134
rect 334928 74866 335248 74898
rect 340094 74550 340154 85443
rect 340094 74490 340522 74550
rect 340091 73540 340157 73541
rect 340091 73476 340092 73540
rect 340156 73476 340157 73540
rect 340091 73475 340157 73476
rect 340094 69730 340154 73475
rect 339542 69670 340154 69730
rect 339542 59941 339602 69670
rect 340462 68370 340522 74490
rect 340094 68310 340522 68370
rect 339539 59940 339605 59941
rect 339539 59876 339540 59940
rect 339604 59876 339605 59940
rect 339539 59875 339605 59876
rect 303294 52954 303914 58000
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 299979 3636 300045 3637
rect 299979 3572 299980 3636
rect 300044 3572 300045 3636
rect 299979 3571 300045 3572
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 57454 308414 58000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 25954 312914 58000
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 30454 317414 58000
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 34954 321914 58000
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 43954 330914 58000
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 48454 335414 58000
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 52954 339914 58000
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 340094 3501 340154 68310
rect 340830 4861 340890 108291
rect 342299 106180 342365 106181
rect 342299 106116 342300 106180
rect 342364 106116 342365 106180
rect 342299 106115 342365 106116
rect 341011 95300 341077 95301
rect 341011 95236 341012 95300
rect 341076 95236 341077 95300
rect 341011 95235 341077 95236
rect 341014 60213 341074 95235
rect 342302 85509 342362 106115
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 342299 85508 342365 85509
rect 342299 85444 342300 85508
rect 342364 85444 342365 85508
rect 342299 85443 342365 85444
rect 342483 84420 342549 84421
rect 342483 84356 342484 84420
rect 342548 84356 342549 84420
rect 342483 84355 342549 84356
rect 342299 82244 342365 82245
rect 342299 82180 342300 82244
rect 342364 82180 342365 82244
rect 342299 82179 342365 82180
rect 341379 79388 341445 79389
rect 341379 79324 341380 79388
rect 341444 79324 341445 79388
rect 341379 79323 341445 79324
rect 341195 71364 341261 71365
rect 341195 71300 341196 71364
rect 341260 71300 341261 71364
rect 341195 71299 341261 71300
rect 341198 61437 341258 71299
rect 341195 61436 341261 61437
rect 341195 61372 341196 61436
rect 341260 61372 341261 61436
rect 341195 61371 341261 61372
rect 341011 60212 341077 60213
rect 341011 60148 341012 60212
rect 341076 60148 341077 60212
rect 341011 60147 341077 60148
rect 340827 4860 340893 4861
rect 340827 4796 340828 4860
rect 340892 4796 340893 4860
rect 340827 4795 340893 4796
rect 340091 3500 340157 3501
rect 340091 3436 340092 3500
rect 340156 3436 340157 3500
rect 340091 3435 340157 3436
rect 341382 3365 341442 79323
rect 342302 10437 342362 82179
rect 342486 58581 342546 84355
rect 342667 77892 342733 77893
rect 342667 77828 342668 77892
rect 342732 77828 342733 77892
rect 342667 77827 342733 77828
rect 342670 60077 342730 77827
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 342667 60076 342733 60077
rect 342667 60012 342668 60076
rect 342732 60012 342733 60076
rect 342667 60011 342733 60012
rect 342483 58580 342549 58581
rect 342483 58516 342484 58580
rect 342548 58516 342549 58580
rect 342483 58515 342549 58516
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 342299 10436 342365 10437
rect 342299 10372 342300 10436
rect 342364 10372 342365 10436
rect 342299 10371 342365 10372
rect 341379 3364 341445 3365
rect 341379 3300 341380 3364
rect 341444 3300 341445 3364
rect 341379 3299 341445 3300
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 349110 3637 349170 518875
rect 352794 498454 353414 533898
rect 349659 498268 349725 498269
rect 349659 498204 349660 498268
rect 349724 498204 349725 498268
rect 349659 498203 349725 498204
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 349662 60349 349722 498203
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 332000 353414 353898
rect 351867 320244 351933 320245
rect 351867 320180 351868 320244
rect 351932 320180 351933 320244
rect 351867 320179 351933 320180
rect 351870 276725 351930 320179
rect 351867 276724 351933 276725
rect 351867 276660 351868 276724
rect 351932 276660 351933 276724
rect 351867 276659 351933 276660
rect 352794 246454 353414 278000
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 349659 60348 349725 60349
rect 349659 60284 349660 60348
rect 349724 60284 349725 60348
rect 349659 60283 349725 60284
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 349107 3636 349173 3637
rect 349107 3572 349108 3636
rect 349172 3572 349173 3636
rect 349107 3571 349173 3572
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 -6106 353414 29898
rect 355182 19413 355242 640323
rect 355366 178125 355426 640459
rect 359043 554300 359109 554301
rect 359043 554236 359044 554300
rect 359108 554236 359109 554300
rect 359043 554235 359109 554236
rect 358859 554028 358925 554029
rect 358859 553964 358860 554028
rect 358924 553964 358925 554028
rect 358859 553963 358925 553964
rect 358307 553484 358373 553485
rect 358307 553420 358308 553484
rect 358372 553420 358373 553484
rect 358307 553419 358373 553420
rect 358123 550628 358189 550629
rect 358123 550564 358124 550628
rect 358188 550564 358189 550628
rect 358123 550563 358189 550564
rect 358126 540701 358186 550563
rect 358310 547093 358370 553419
rect 358675 551988 358741 551989
rect 358675 551924 358676 551988
rect 358740 551924 358741 551988
rect 358675 551923 358741 551924
rect 358491 551852 358557 551853
rect 358491 551788 358492 551852
rect 358556 551788 358557 551852
rect 358491 551787 358557 551788
rect 358307 547092 358373 547093
rect 358307 547028 358308 547092
rect 358372 547028 358373 547092
rect 358307 547027 358373 547028
rect 358123 540700 358189 540701
rect 358123 540636 358124 540700
rect 358188 540636 358189 540700
rect 358123 540635 358189 540636
rect 358494 530637 358554 551787
rect 358491 530636 358557 530637
rect 358491 530572 358492 530636
rect 358556 530572 358557 530636
rect 358491 530571 358557 530572
rect 358678 502349 358738 551923
rect 358862 505069 358922 553963
rect 359046 541109 359106 554235
rect 359043 541108 359109 541109
rect 359043 541044 359044 541108
rect 359108 541044 359109 541108
rect 359043 541043 359109 541044
rect 358859 505068 358925 505069
rect 358859 505004 358860 505068
rect 358924 505004 358925 505068
rect 358859 505003 358925 505004
rect 358675 502348 358741 502349
rect 358675 502284 358676 502348
rect 358740 502284 358741 502348
rect 358675 502283 358741 502284
rect 359414 501261 359474 642091
rect 361794 642000 362414 650898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 642000 366914 655398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 642000 371414 659898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 642000 375914 664398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 642000 380414 668898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 642000 384914 673398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642361 389414 677898
rect 388794 642125 388826 642361
rect 389062 642125 389146 642361
rect 389382 642125 389414 642361
rect 388794 642000 389414 642125
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 642000 393914 646398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 401547 661332 401613 661333
rect 401547 661268 401548 661332
rect 401612 661268 401613 661332
rect 401547 661267 401613 661268
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 642000 398414 650898
rect 398603 642020 398669 642021
rect 398603 641956 398604 642020
rect 398668 641956 398669 642020
rect 398603 641955 398669 641956
rect 363459 641748 363525 641749
rect 363459 641684 363460 641748
rect 363524 641684 363525 641748
rect 363459 641683 363525 641684
rect 362539 639980 362605 639981
rect 362539 639916 362540 639980
rect 362604 639916 362605 639980
rect 362539 639915 362605 639916
rect 362355 639572 362421 639573
rect 362355 639508 362356 639572
rect 362420 639508 362421 639572
rect 362355 639507 362421 639508
rect 360699 598364 360765 598365
rect 360699 598300 360700 598364
rect 360764 598300 360765 598364
rect 360699 598299 360765 598300
rect 360702 528570 360762 598299
rect 362358 569261 362418 639507
rect 362542 596869 362602 639915
rect 362723 639436 362789 639437
rect 362723 639372 362724 639436
rect 362788 639372 362789 639436
rect 362723 639371 362789 639372
rect 362539 596868 362605 596869
rect 362539 596804 362540 596868
rect 362604 596804 362605 596868
rect 362539 596803 362605 596804
rect 362539 583132 362605 583133
rect 362539 583068 362540 583132
rect 362604 583068 362605 583132
rect 362539 583067 362605 583068
rect 362355 569260 362421 569261
rect 362355 569196 362356 569260
rect 362420 569196 362421 569260
rect 362355 569195 362421 569196
rect 361619 565180 361685 565181
rect 361619 565116 361620 565180
rect 361684 565116 361685 565180
rect 361619 565115 361685 565116
rect 361435 563956 361501 563957
rect 361435 563892 361436 563956
rect 361500 563892 361501 563956
rect 361435 563891 361501 563892
rect 360518 528510 360762 528570
rect 360518 526965 360578 528510
rect 360515 526964 360581 526965
rect 360515 526900 360516 526964
rect 360580 526900 360581 526964
rect 360515 526899 360581 526900
rect 359411 501260 359477 501261
rect 359411 501196 359412 501260
rect 359476 501196 359477 501260
rect 359411 501195 359477 501196
rect 361438 499901 361498 563891
rect 361622 499901 361682 565115
rect 361435 499900 361501 499901
rect 361435 499836 361436 499900
rect 361500 499836 361501 499900
rect 361435 499835 361501 499836
rect 361619 499900 361685 499901
rect 361619 499836 361620 499900
rect 361684 499836 361685 499900
rect 361619 499835 361685 499836
rect 362542 498133 362602 583067
rect 362726 561101 362786 639371
rect 362723 561100 362789 561101
rect 362723 561036 362724 561100
rect 362788 561036 362789 561100
rect 362723 561035 362789 561036
rect 362907 560284 362973 560285
rect 362907 560220 362908 560284
rect 362972 560220 362973 560284
rect 362907 560219 362973 560220
rect 362539 498132 362605 498133
rect 362539 498068 362540 498132
rect 362604 498068 362605 498132
rect 362539 498067 362605 498068
rect 357294 466954 357914 498000
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 355363 178124 355429 178125
rect 355363 178060 355364 178124
rect 355428 178060 355429 178124
rect 355363 178059 355429 178060
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 355179 19412 355245 19413
rect 355179 19348 355180 19412
rect 355244 19348 355245 19412
rect 355179 19347 355245 19348
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 471454 362414 498000
rect 362910 497861 362970 560219
rect 363462 558925 363522 641683
rect 364011 639436 364077 639437
rect 364011 639372 364012 639436
rect 364076 639372 364077 639436
rect 364011 639371 364077 639372
rect 364014 585717 364074 639371
rect 379568 619954 379888 619986
rect 379568 619718 379610 619954
rect 379846 619718 379888 619954
rect 379568 619634 379888 619718
rect 379568 619398 379610 619634
rect 379846 619398 379888 619634
rect 379568 619366 379888 619398
rect 364208 615454 364528 615486
rect 364208 615218 364250 615454
rect 364486 615218 364528 615454
rect 364208 615134 364528 615218
rect 364208 614898 364250 615134
rect 364486 614898 364528 615134
rect 364208 614866 364528 614898
rect 394928 615454 395248 615486
rect 394928 615218 394970 615454
rect 395206 615218 395248 615454
rect 394928 615134 395248 615218
rect 394928 614898 394970 615134
rect 395206 614898 395248 615134
rect 394928 614866 395248 614898
rect 366219 598228 366285 598229
rect 366219 598164 366220 598228
rect 366284 598164 366285 598228
rect 366219 598163 366285 598164
rect 369899 598228 369965 598229
rect 369899 598164 369900 598228
rect 369964 598164 369965 598228
rect 369899 598163 369965 598164
rect 379283 598228 379349 598229
rect 379283 598164 379284 598228
rect 379348 598164 379349 598228
rect 379283 598163 379349 598164
rect 364011 585716 364077 585717
rect 364011 585652 364012 585716
rect 364076 585652 364077 585716
rect 364011 585651 364077 585652
rect 364747 560964 364813 560965
rect 364747 560900 364748 560964
rect 364812 560900 364813 560964
rect 364747 560899 364813 560900
rect 363459 558924 363525 558925
rect 363459 558860 363460 558924
rect 363524 558860 363525 558924
rect 363459 558859 363525 558860
rect 364208 543454 364528 543486
rect 364208 543218 364250 543454
rect 364486 543218 364528 543454
rect 364208 543134 364528 543218
rect 364208 542898 364250 543134
rect 364486 542898 364528 543134
rect 364208 542866 364528 542898
rect 364208 507454 364528 507486
rect 364208 507218 364250 507454
rect 364486 507218 364528 507454
rect 364208 507134 364528 507218
rect 364208 506898 364250 507134
rect 364486 506898 364528 507134
rect 364208 506866 364528 506898
rect 364750 499901 364810 560899
rect 364747 499900 364813 499901
rect 364747 499836 364748 499900
rect 364812 499836 364813 499900
rect 364747 499835 364813 499836
rect 366222 499493 366282 598163
rect 368243 581772 368309 581773
rect 368243 581708 368244 581772
rect 368308 581708 368309 581772
rect 368243 581707 368309 581708
rect 368246 499901 368306 581707
rect 368427 568036 368493 568037
rect 368427 567972 368428 568036
rect 368492 567972 368493 568036
rect 368427 567971 368493 567972
rect 368430 518910 368490 567971
rect 368430 518850 368674 518910
rect 368614 499901 368674 518850
rect 368243 499900 368309 499901
rect 368243 499836 368244 499900
rect 368308 499836 368309 499900
rect 368243 499835 368309 499836
rect 368611 499900 368677 499901
rect 368611 499836 368612 499900
rect 368676 499836 368677 499900
rect 368611 499835 368677 499836
rect 366219 499492 366285 499493
rect 366219 499428 366220 499492
rect 366284 499428 366285 499492
rect 366219 499427 366285 499428
rect 369902 498949 369962 598163
rect 370794 588454 371414 598000
rect 373211 597684 373277 597685
rect 373211 597620 373212 597684
rect 373276 597620 373277 597684
rect 373211 597619 373277 597620
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370083 571980 370149 571981
rect 370083 571916 370084 571980
rect 370148 571916 370149 571980
rect 370083 571915 370149 571916
rect 370086 499901 370146 571915
rect 370794 552361 371414 587898
rect 371739 580412 371805 580413
rect 371739 580348 371740 580412
rect 371804 580348 371805 580412
rect 371739 580347 371805 580348
rect 370794 552125 370826 552361
rect 371062 552125 371146 552361
rect 371382 552125 371414 552361
rect 370794 552000 371414 552125
rect 370083 499900 370149 499901
rect 370083 499836 370084 499900
rect 370148 499836 370149 499900
rect 370083 499835 370149 499836
rect 369899 498948 369965 498949
rect 369899 498884 369900 498948
rect 369964 498884 369965 498948
rect 369899 498883 369965 498884
rect 362907 497860 362973 497861
rect 362907 497796 362908 497860
rect 362972 497796 362973 497860
rect 362907 497795 362973 497796
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 475954 366914 498000
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 480454 371414 498000
rect 371742 497997 371802 580347
rect 373214 499493 373274 597619
rect 375294 592954 375914 598000
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 373395 592652 373461 592653
rect 373395 592588 373396 592652
rect 373460 592588 373461 592652
rect 373395 592587 373461 592588
rect 375294 592634 375914 592718
rect 373211 499492 373277 499493
rect 373211 499428 373212 499492
rect 373276 499428 373277 499492
rect 373211 499427 373277 499428
rect 371739 497996 371805 497997
rect 371739 497932 371740 497996
rect 371804 497932 371805 497996
rect 371739 497931 371805 497932
rect 373398 497317 373458 592587
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 373763 565044 373829 565045
rect 373763 564980 373764 565044
rect 373828 564980 373829 565044
rect 373763 564979 373829 564980
rect 373766 499901 373826 564979
rect 375294 556954 375914 592398
rect 376155 580276 376221 580277
rect 376155 580212 376156 580276
rect 376220 580212 376221 580276
rect 376155 580211 376221 580212
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 552000 375914 556398
rect 373763 499900 373829 499901
rect 373763 499836 373764 499900
rect 373828 499836 373829 499900
rect 373763 499835 373829 499836
rect 376158 499493 376218 580211
rect 376891 568172 376957 568173
rect 376891 568108 376892 568172
rect 376956 568108 376957 568172
rect 376891 568107 376957 568108
rect 376339 568036 376405 568037
rect 376339 567972 376340 568036
rect 376404 567972 376405 568036
rect 376339 567971 376405 567972
rect 376342 499901 376402 567971
rect 376894 499901 376954 568107
rect 376339 499900 376405 499901
rect 376339 499836 376340 499900
rect 376404 499836 376405 499900
rect 376339 499835 376405 499836
rect 376891 499900 376957 499901
rect 376891 499836 376892 499900
rect 376956 499836 376957 499900
rect 376891 499835 376957 499836
rect 376155 499492 376221 499493
rect 376155 499428 376156 499492
rect 376220 499428 376221 499492
rect 376155 499427 376221 499428
rect 373395 497316 373461 497317
rect 373395 497252 373396 497316
rect 373460 497252 373461 497316
rect 373395 497251 373461 497252
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 484954 375914 498000
rect 379286 497997 379346 598163
rect 379794 597454 380414 598000
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 382779 595508 382845 595509
rect 382779 595444 382780 595508
rect 382844 595444 382845 595508
rect 382779 595443 382845 595444
rect 380939 581636 381005 581637
rect 380939 581572 380940 581636
rect 381004 581572 381005 581636
rect 380939 581571 381005 581572
rect 380571 566404 380637 566405
rect 380571 566340 380572 566404
rect 380636 566340 380637 566404
rect 380571 566339 380637 566340
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 552000 380414 560898
rect 379568 511954 379888 511986
rect 379568 511718 379610 511954
rect 379846 511718 379888 511954
rect 379568 511634 379888 511718
rect 379568 511398 379610 511634
rect 379846 511398 379888 511634
rect 379568 511366 379888 511398
rect 380574 499901 380634 566339
rect 380942 499901 381002 581571
rect 382782 499901 382842 595443
rect 392531 586396 392597 586397
rect 392531 586332 392532 586396
rect 392596 586332 392597 586396
rect 392531 586331 392597 586332
rect 387011 583812 387077 583813
rect 387011 583748 387012 583812
rect 387076 583748 387077 583812
rect 387011 583747 387077 583748
rect 384067 576876 384133 576877
rect 384067 576812 384068 576876
rect 384132 576812 384133 576876
rect 384067 576811 384133 576812
rect 380571 499900 380637 499901
rect 380571 499836 380572 499900
rect 380636 499836 380637 499900
rect 380571 499835 380637 499836
rect 380939 499900 381005 499901
rect 380939 499836 380940 499900
rect 381004 499836 381005 499900
rect 380939 499835 381005 499836
rect 382779 499900 382845 499901
rect 382779 499836 382780 499900
rect 382844 499836 382845 499900
rect 382779 499835 382845 499836
rect 384070 498133 384130 576811
rect 385539 560284 385605 560285
rect 385539 560220 385540 560284
rect 385604 560220 385605 560284
rect 385539 560219 385605 560220
rect 385542 499901 385602 560219
rect 385539 499900 385605 499901
rect 385539 499836 385540 499900
rect 385604 499836 385605 499900
rect 385539 499835 385605 499836
rect 384067 498132 384133 498133
rect 384067 498068 384068 498132
rect 384132 498068 384133 498132
rect 384067 498067 384133 498068
rect 379283 497996 379349 497997
rect 379283 497932 379284 497996
rect 379348 497932 379349 497996
rect 379283 497931 379349 497932
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 489454 380414 498000
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 493954 384914 498000
rect 387014 497725 387074 583747
rect 388299 582996 388365 582997
rect 388299 582932 388300 582996
rect 388364 582932 388365 582996
rect 388299 582931 388365 582932
rect 388302 498133 388362 582931
rect 391979 581908 392045 581909
rect 391979 581844 391980 581908
rect 392044 581844 392045 581908
rect 391979 581843 392045 581844
rect 391059 574836 391125 574837
rect 391059 574772 391060 574836
rect 391124 574772 391125 574836
rect 391059 574771 391125 574772
rect 389587 574700 389653 574701
rect 389587 574636 389588 574700
rect 389652 574636 389653 574700
rect 389587 574635 389653 574636
rect 389590 499901 389650 574635
rect 389587 499900 389653 499901
rect 389587 499836 389588 499900
rect 389652 499836 389653 499900
rect 389587 499835 389653 499836
rect 391062 499629 391122 574771
rect 391982 499901 392042 581843
rect 391979 499900 392045 499901
rect 391979 499836 391980 499900
rect 392044 499836 392045 499900
rect 391979 499835 392045 499836
rect 392534 499765 392594 586331
rect 396579 573340 396645 573341
rect 396579 573276 396580 573340
rect 396644 573276 396645 573340
rect 396579 573275 396645 573276
rect 394928 543454 395248 543486
rect 394928 543218 394970 543454
rect 395206 543218 395248 543454
rect 394928 543134 395248 543218
rect 394928 542898 394970 543134
rect 395206 542898 395248 543134
rect 394928 542866 395248 542898
rect 394928 507454 395248 507486
rect 394928 507218 394970 507454
rect 395206 507218 395248 507454
rect 394928 507134 395248 507218
rect 394928 506898 394970 507134
rect 395206 506898 395248 507134
rect 394928 506866 395248 506898
rect 396582 499901 396642 573275
rect 398606 539610 398666 641955
rect 400259 563820 400325 563821
rect 400259 563756 400260 563820
rect 400324 563756 400325 563820
rect 400259 563755 400325 563756
rect 398787 563684 398853 563685
rect 398787 563620 398788 563684
rect 398852 563620 398853 563684
rect 398787 563619 398853 563620
rect 398238 539550 398666 539610
rect 398238 532130 398298 539550
rect 398790 537570 398850 563619
rect 399155 562324 399221 562325
rect 399155 562260 399156 562324
rect 399220 562260 399221 562324
rect 399155 562259 399221 562260
rect 398971 551308 399037 551309
rect 398971 551244 398972 551308
rect 399036 551244 399037 551308
rect 398971 551243 399037 551244
rect 398974 538230 399034 551243
rect 399158 539610 399218 562259
rect 399339 550628 399405 550629
rect 399339 550564 399340 550628
rect 399404 550564 399405 550628
rect 399339 550563 399405 550564
rect 399342 543829 399402 550563
rect 399339 543828 399405 543829
rect 399339 543764 399340 543828
rect 399404 543764 399405 543828
rect 399339 543763 399405 543764
rect 399158 539550 399954 539610
rect 398974 538170 399402 538230
rect 398422 537510 398850 537570
rect 398422 535530 398482 537510
rect 399342 535669 399402 538170
rect 399339 535668 399405 535669
rect 399339 535604 399340 535668
rect 399404 535604 399405 535668
rect 399339 535603 399405 535604
rect 398422 535470 399218 535530
rect 399158 534850 399218 535470
rect 399158 534790 399770 534850
rect 399339 533220 399405 533221
rect 399339 533156 399340 533220
rect 399404 533156 399405 533220
rect 399339 533155 399405 533156
rect 399342 532810 399402 533155
rect 398974 532750 399402 532810
rect 398238 532070 398666 532130
rect 396579 499900 396645 499901
rect 396579 499836 396580 499900
rect 396644 499836 396645 499900
rect 396579 499835 396645 499836
rect 398606 499765 398666 532070
rect 398974 514770 399034 532750
rect 399710 531450 399770 534790
rect 399158 531390 399770 531450
rect 399158 521250 399218 531390
rect 399894 529950 399954 539550
rect 399342 529890 399954 529950
rect 399342 521661 399402 529890
rect 399339 521660 399405 521661
rect 399339 521596 399340 521660
rect 399404 521596 399405 521660
rect 399339 521595 399405 521596
rect 399158 521190 399402 521250
rect 399342 518805 399402 521190
rect 399339 518804 399405 518805
rect 399339 518740 399340 518804
rect 399404 518740 399405 518804
rect 399339 518739 399405 518740
rect 398974 514710 399402 514770
rect 399342 507789 399402 514710
rect 399339 507788 399405 507789
rect 399339 507724 399340 507788
rect 399404 507724 399405 507788
rect 399339 507723 399405 507724
rect 400262 501465 400322 563755
rect 400443 558244 400509 558245
rect 400443 558180 400444 558244
rect 400508 558180 400509 558244
rect 400443 558179 400509 558180
rect 400446 504865 400506 558179
rect 400627 554164 400693 554165
rect 400627 554100 400628 554164
rect 400692 554100 400693 554164
rect 400627 554099 400693 554100
rect 400630 537845 400690 554099
rect 400811 551444 400877 551445
rect 400811 551380 400812 551444
rect 400876 551380 400877 551444
rect 400811 551379 400877 551380
rect 400814 547773 400874 551379
rect 401550 549269 401610 661267
rect 402294 655954 402914 691398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 403019 662828 403085 662829
rect 403019 662764 403020 662828
rect 403084 662764 403085 662828
rect 403019 662763 403085 662764
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 642000 402914 655398
rect 401731 555388 401797 555389
rect 401731 555324 401732 555388
rect 401796 555324 401797 555388
rect 401731 555323 401797 555324
rect 401547 549268 401613 549269
rect 401547 549204 401548 549268
rect 401612 549204 401613 549268
rect 401547 549203 401613 549204
rect 400811 547772 400877 547773
rect 400811 547708 400812 547772
rect 400876 547708 400877 547772
rect 400811 547707 400877 547708
rect 400627 537844 400693 537845
rect 400627 537780 400628 537844
rect 400692 537780 400693 537844
rect 400627 537779 400693 537780
rect 401734 508333 401794 555323
rect 403022 539613 403082 662763
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 404859 596868 404925 596869
rect 404859 596804 404860 596868
rect 404924 596804 404925 596868
rect 404859 596803 404925 596804
rect 403571 552124 403637 552125
rect 403571 552060 403572 552124
rect 403636 552060 403637 552124
rect 403571 552059 403637 552060
rect 403019 539612 403085 539613
rect 403019 539548 403020 539612
rect 403084 539548 403085 539612
rect 403019 539547 403085 539548
rect 401731 508332 401797 508333
rect 401731 508268 401732 508332
rect 401796 508268 401797 508332
rect 401731 508267 401797 508268
rect 400443 504864 400509 504865
rect 400443 504800 400444 504864
rect 400508 504800 400509 504864
rect 400443 504799 400509 504800
rect 400259 501464 400325 501465
rect 400259 501400 400260 501464
rect 400324 501400 400325 501464
rect 400259 501399 400325 501400
rect 392531 499764 392597 499765
rect 392531 499700 392532 499764
rect 392596 499700 392597 499764
rect 392531 499699 392597 499700
rect 398603 499764 398669 499765
rect 398603 499700 398604 499764
rect 398668 499700 398669 499764
rect 398603 499699 398669 499700
rect 391059 499628 391125 499629
rect 391059 499564 391060 499628
rect 391124 499564 391125 499628
rect 391059 499563 391125 499564
rect 388299 498132 388365 498133
rect 388299 498068 388300 498132
rect 388364 498068 388365 498132
rect 388299 498067 388365 498068
rect 387011 497724 387077 497725
rect 387011 497660 387012 497724
rect 387076 497660 387077 497724
rect 387011 497659 387077 497660
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 462454 389414 498000
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 466954 393914 498000
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 471454 398414 498000
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 475954 402914 498000
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 403574 177309 403634 552059
rect 404862 509421 404922 596803
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 404859 509420 404925 509421
rect 404859 509356 404860 509420
rect 404924 509356 404925 509420
rect 404859 509355 404925 509356
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 403571 177308 403637 177309
rect 403571 177244 403572 177308
rect 403636 177244 403637 177308
rect 403571 177243 403637 177244
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 481587 662692 481653 662693
rect 481587 662628 481588 662692
rect 481652 662628 481653 662692
rect 481587 662627 481653 662628
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 642000 479414 659898
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 478794 588454 479414 598000
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 532000 479414 551898
rect 481590 532677 481650 662627
rect 483294 642000 483914 664398
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 484899 661060 484965 661061
rect 484899 660996 484900 661060
rect 484964 660996 484965 661060
rect 484899 660995 484965 660996
rect 484208 615454 484528 615486
rect 484208 615218 484250 615454
rect 484486 615218 484528 615454
rect 484208 615134 484528 615218
rect 484208 614898 484250 615134
rect 484486 614898 484528 615134
rect 484208 614866 484528 614898
rect 483294 592954 483914 598000
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 481587 532676 481653 532677
rect 481587 532612 481588 532676
rect 481652 532612 481653 532676
rect 481587 532611 481653 532612
rect 483294 532000 483914 556398
rect 484902 532677 484962 660995
rect 487794 642000 488414 668898
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 489131 660244 489197 660245
rect 489131 660180 489132 660244
rect 489196 660180 489197 660244
rect 489131 660179 489197 660180
rect 487794 597454 488414 598000
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 484899 532676 484965 532677
rect 484899 532612 484900 532676
rect 484964 532612 484965 532676
rect 484899 532611 484965 532612
rect 487794 532000 488414 560898
rect 489134 532677 489194 660179
rect 492294 642000 492914 673398
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 495387 662556 495453 662557
rect 495387 662492 495388 662556
rect 495452 662492 495453 662556
rect 495387 662491 495453 662492
rect 489131 532676 489197 532677
rect 489131 532612 489132 532676
rect 489196 532612 489197 532676
rect 489131 532611 489197 532612
rect 484163 529956 484229 529957
rect 484163 529892 484164 529956
rect 484228 529892 484229 529956
rect 484163 529891 484229 529892
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 480454 479414 498000
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 484954 483914 498000
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 484166 4045 484226 529891
rect 489683 529548 489749 529549
rect 489683 529484 489684 529548
rect 489748 529484 489749 529548
rect 489683 529483 489749 529484
rect 487892 511954 488212 511986
rect 487892 511718 487934 511954
rect 488170 511718 488212 511954
rect 487892 511634 488212 511718
rect 487892 511398 487934 511634
rect 488170 511398 488212 511634
rect 487892 511366 488212 511398
rect 484418 507454 484738 507486
rect 484418 507218 484460 507454
rect 484696 507218 484738 507454
rect 484418 507134 484738 507218
rect 484418 506898 484460 507134
rect 484696 506898 484738 507134
rect 484418 506866 484738 506898
rect 487794 489454 488414 498000
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 489686 39269 489746 529483
rect 494840 511954 495160 511986
rect 494840 511718 494882 511954
rect 495118 511718 495160 511954
rect 494840 511634 495160 511718
rect 494840 511398 494882 511634
rect 495118 511398 495160 511634
rect 494840 511366 495160 511398
rect 491366 507454 491686 507486
rect 491366 507218 491408 507454
rect 491644 507218 491686 507454
rect 491366 507134 491686 507218
rect 491366 506898 491408 507134
rect 491644 506898 491686 507134
rect 491366 506866 491686 506898
rect 495390 499901 495450 662491
rect 496794 642361 497414 677898
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 499435 661060 499501 661061
rect 499435 660996 499436 661060
rect 499500 660996 499501 661060
rect 499435 660995 499501 660996
rect 496794 642125 496826 642361
rect 497062 642125 497146 642361
rect 497382 642125 497414 642361
rect 496794 642000 497414 642125
rect 496794 570454 497414 598000
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 532000 497414 533898
rect 499438 532541 499498 660995
rect 501294 646954 501914 682398
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 502011 659836 502077 659837
rect 502011 659772 502012 659836
rect 502076 659772 502077 659836
rect 502011 659771 502077 659772
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 642000 501914 646398
rect 499568 619954 499888 619986
rect 499568 619718 499610 619954
rect 499846 619718 499888 619954
rect 499568 619634 499888 619718
rect 499568 619398 499610 619634
rect 499846 619398 499888 619634
rect 499568 619366 499888 619398
rect 501294 574954 501914 598000
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 499435 532540 499501 532541
rect 499435 532476 499436 532540
rect 499500 532476 499501 532540
rect 499435 532475 499501 532476
rect 501294 532000 501914 538398
rect 502014 532677 502074 659771
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 642000 506414 650898
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 512131 661196 512197 661197
rect 512131 661132 512132 661196
rect 512196 661132 512197 661196
rect 512131 661131 512197 661132
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 642000 510914 655398
rect 505794 579454 506414 598000
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 502011 532676 502077 532677
rect 502011 532612 502012 532676
rect 502076 532612 502077 532676
rect 502011 532611 502077 532612
rect 505794 532000 506414 542898
rect 510294 583954 510914 598000
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 532000 510914 547398
rect 502379 529548 502445 529549
rect 502379 529484 502380 529548
rect 502444 529484 502445 529548
rect 502379 529483 502445 529484
rect 503667 529548 503733 529549
rect 503667 529484 503668 529548
rect 503732 529484 503733 529548
rect 503667 529483 503733 529484
rect 501788 511954 502108 511986
rect 501788 511718 501830 511954
rect 502066 511718 502108 511954
rect 501788 511634 502108 511718
rect 501788 511398 501830 511634
rect 502066 511398 502108 511634
rect 501788 511366 502108 511398
rect 498314 507454 498634 507486
rect 498314 507218 498356 507454
rect 498592 507218 498634 507454
rect 498314 507134 498634 507218
rect 498314 506898 498356 507134
rect 498592 506898 498634 507134
rect 498314 506866 498634 506898
rect 495387 499900 495453 499901
rect 495387 499836 495388 499900
rect 495452 499836 495453 499900
rect 495387 499835 495453 499836
rect 502382 498813 502442 529483
rect 502379 498812 502445 498813
rect 502379 498748 502380 498812
rect 502444 498748 502445 498812
rect 502379 498747 502445 498748
rect 492294 493954 492914 498000
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 489683 39268 489749 39269
rect 489683 39204 489684 39268
rect 489748 39204 489749 39268
rect 489683 39203 489749 39204
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 484163 4044 484229 4045
rect 484163 3980 484164 4044
rect 484228 3980 484229 4044
rect 484163 3979 484229 3980
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 462454 497414 498000
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 466954 501914 498000
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 503670 8941 503730 529483
rect 509371 527508 509437 527509
rect 509371 527444 509372 527508
rect 509436 527444 509437 527508
rect 509371 527443 509437 527444
rect 509374 521670 509434 527443
rect 509006 521610 509434 521670
rect 505262 507454 505582 507486
rect 505262 507218 505304 507454
rect 505540 507218 505582 507454
rect 505262 507134 505582 507218
rect 505262 506898 505304 507134
rect 505540 506898 505582 507134
rect 505262 506866 505582 506898
rect 505794 471454 506414 498000
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 503667 8940 503733 8941
rect 503667 8876 503668 8940
rect 503732 8876 503733 8940
rect 503667 8875 503733 8876
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 3454 506414 38898
rect 509006 10301 509066 521610
rect 512134 512821 512194 661131
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 642000 515414 659898
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 642000 519914 664398
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 642000 524414 668898
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 514928 615454 515248 615486
rect 514928 615218 514970 615454
rect 515206 615218 515248 615454
rect 514928 615134 515248 615218
rect 514928 614898 514970 615134
rect 515206 614898 515248 615134
rect 514928 614866 515248 614898
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 514794 588454 515414 598000
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 512131 512820 512197 512821
rect 512131 512756 512132 512820
rect 512196 512756 512197 512820
rect 512131 512755 512197 512756
rect 510294 475954 510914 498000
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 509003 10300 509069 10301
rect 509003 10236 509004 10300
rect 509068 10236 509069 10300
rect 509003 10235 509069 10236
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 592954 519914 598000
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 597454 524414 598000
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 71610 655718 71846 655954
rect 71610 655398 71846 655634
rect 102330 655718 102566 655954
rect 102330 655398 102566 655634
rect 133050 655718 133286 655954
rect 133050 655398 133286 655634
rect 163770 655718 164006 655954
rect 163770 655398 164006 655634
rect 194490 655718 194726 655954
rect 194490 655398 194726 655634
rect 225210 655718 225446 655954
rect 225210 655398 225446 655634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 56250 651218 56486 651454
rect 56250 650898 56486 651134
rect 86970 651218 87206 651454
rect 86970 650898 87206 651134
rect 117690 651218 117926 651454
rect 117690 650898 117926 651134
rect 148410 651218 148646 651454
rect 148410 650898 148646 651134
rect 179130 651218 179366 651454
rect 179130 650898 179366 651134
rect 209850 651218 210086 651454
rect 209850 650898 210086 651134
rect 240570 651218 240806 651454
rect 240570 650898 240806 651134
rect 71610 619718 71846 619954
rect 71610 619398 71846 619634
rect 102330 619718 102566 619954
rect 102330 619398 102566 619634
rect 133050 619718 133286 619954
rect 133050 619398 133286 619634
rect 163770 619718 164006 619954
rect 163770 619398 164006 619634
rect 194490 619718 194726 619954
rect 194490 619398 194726 619634
rect 225210 619718 225446 619954
rect 225210 619398 225446 619634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 56250 615218 56486 615454
rect 56250 614898 56486 615134
rect 86970 615218 87206 615454
rect 86970 614898 87206 615134
rect 117690 615218 117926 615454
rect 117690 614898 117926 615134
rect 148410 615218 148646 615454
rect 148410 614898 148646 615134
rect 179130 615218 179366 615454
rect 179130 614898 179366 615134
rect 209850 615218 210086 615454
rect 209850 614898 210086 615134
rect 240570 615218 240806 615454
rect 240570 614898 240806 615134
rect 71610 583718 71846 583954
rect 71610 583398 71846 583634
rect 102330 583718 102566 583954
rect 102330 583398 102566 583634
rect 133050 583718 133286 583954
rect 133050 583398 133286 583634
rect 163770 583718 164006 583954
rect 163770 583398 164006 583634
rect 194490 583718 194726 583954
rect 194490 583398 194726 583634
rect 225210 583718 225446 583954
rect 225210 583398 225446 583634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 56250 579218 56486 579454
rect 56250 578898 56486 579134
rect 86970 579218 87206 579454
rect 86970 578898 87206 579134
rect 117690 579218 117926 579454
rect 117690 578898 117926 579134
rect 148410 579218 148646 579454
rect 148410 578898 148646 579134
rect 179130 579218 179366 579454
rect 179130 578898 179366 579134
rect 209850 579218 210086 579454
rect 209850 578898 210086 579134
rect 240570 579218 240806 579454
rect 240570 578898 240806 579134
rect 71610 547718 71846 547954
rect 71610 547398 71846 547634
rect 102330 547718 102566 547954
rect 102330 547398 102566 547634
rect 133050 547718 133286 547954
rect 133050 547398 133286 547634
rect 163770 547718 164006 547954
rect 163770 547398 164006 547634
rect 194490 547718 194726 547954
rect 194490 547398 194726 547634
rect 225210 547718 225446 547954
rect 225210 547398 225446 547634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 56250 543218 56486 543454
rect 56250 542898 56486 543134
rect 86970 543218 87206 543454
rect 86970 542898 87206 543134
rect 117690 543218 117926 543454
rect 117690 542898 117926 543134
rect 148410 543218 148646 543454
rect 148410 542898 148646 543134
rect 179130 543218 179366 543454
rect 179130 542898 179366 543134
rect 209850 543218 210086 543454
rect 209850 542898 210086 543134
rect 240570 543218 240806 543454
rect 240570 542898 240806 543134
rect 71610 511718 71846 511954
rect 71610 511398 71846 511634
rect 102330 511718 102566 511954
rect 102330 511398 102566 511634
rect 133050 511718 133286 511954
rect 133050 511398 133286 511634
rect 163770 511718 164006 511954
rect 163770 511398 164006 511634
rect 194490 511718 194726 511954
rect 194490 511398 194726 511634
rect 225210 511718 225446 511954
rect 225210 511398 225446 511634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 56250 507218 56486 507454
rect 56250 506898 56486 507134
rect 86970 507218 87206 507454
rect 86970 506898 87206 507134
rect 117690 507218 117926 507454
rect 117690 506898 117926 507134
rect 148410 507218 148646 507454
rect 148410 506898 148646 507134
rect 179130 507218 179366 507454
rect 179130 506898 179366 507134
rect 209850 507218 210086 507454
rect 209850 506898 210086 507134
rect 240570 507218 240806 507454
rect 240570 506898 240806 507134
rect 71610 475718 71846 475954
rect 71610 475398 71846 475634
rect 102330 475718 102566 475954
rect 102330 475398 102566 475634
rect 133050 475718 133286 475954
rect 133050 475398 133286 475634
rect 163770 475718 164006 475954
rect 163770 475398 164006 475634
rect 194490 475718 194726 475954
rect 194490 475398 194726 475634
rect 225210 475718 225446 475954
rect 225210 475398 225446 475634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 56250 471218 56486 471454
rect 56250 470898 56486 471134
rect 86970 471218 87206 471454
rect 86970 470898 87206 471134
rect 117690 471218 117926 471454
rect 117690 470898 117926 471134
rect 148410 471218 148646 471454
rect 148410 470898 148646 471134
rect 179130 471218 179366 471454
rect 179130 470898 179366 471134
rect 209850 471218 210086 471454
rect 209850 470898 210086 471134
rect 240570 471218 240806 471454
rect 240570 470898 240806 471134
rect 71610 439718 71846 439954
rect 71610 439398 71846 439634
rect 102330 439718 102566 439954
rect 102330 439398 102566 439634
rect 133050 439718 133286 439954
rect 133050 439398 133286 439634
rect 163770 439718 164006 439954
rect 163770 439398 164006 439634
rect 194490 439718 194726 439954
rect 194490 439398 194726 439634
rect 225210 439718 225446 439954
rect 225210 439398 225446 439634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 56250 435218 56486 435454
rect 56250 434898 56486 435134
rect 86970 435218 87206 435454
rect 86970 434898 87206 435134
rect 117690 435218 117926 435454
rect 117690 434898 117926 435134
rect 148410 435218 148646 435454
rect 148410 434898 148646 435134
rect 179130 435218 179366 435454
rect 179130 434898 179366 435134
rect 209850 435218 210086 435454
rect 209850 434898 210086 435134
rect 240570 435218 240806 435454
rect 240570 434898 240806 435134
rect 71610 403718 71846 403954
rect 71610 403398 71846 403634
rect 102330 403718 102566 403954
rect 102330 403398 102566 403634
rect 133050 403718 133286 403954
rect 133050 403398 133286 403634
rect 163770 403718 164006 403954
rect 163770 403398 164006 403634
rect 194490 403718 194726 403954
rect 194490 403398 194726 403634
rect 225210 403718 225446 403954
rect 225210 403398 225446 403634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 56250 399218 56486 399454
rect 56250 398898 56486 399134
rect 86970 399218 87206 399454
rect 86970 398898 87206 399134
rect 117690 399218 117926 399454
rect 117690 398898 117926 399134
rect 148410 399218 148646 399454
rect 148410 398898 148646 399134
rect 179130 399218 179366 399454
rect 179130 398898 179366 399134
rect 209850 399218 210086 399454
rect 209850 398898 210086 399134
rect 240570 399218 240806 399454
rect 240570 398898 240806 399134
rect 71610 367718 71846 367954
rect 71610 367398 71846 367634
rect 102330 367718 102566 367954
rect 102330 367398 102566 367634
rect 133050 367718 133286 367954
rect 133050 367398 133286 367634
rect 163770 367718 164006 367954
rect 163770 367398 164006 367634
rect 194490 367718 194726 367954
rect 194490 367398 194726 367634
rect 225210 367718 225446 367954
rect 225210 367398 225446 367634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 56250 363218 56486 363454
rect 56250 362898 56486 363134
rect 86970 363218 87206 363454
rect 86970 362898 87206 363134
rect 117690 363218 117926 363454
rect 117690 362898 117926 363134
rect 148410 363218 148646 363454
rect 148410 362898 148646 363134
rect 179130 363218 179366 363454
rect 179130 362898 179366 363134
rect 209850 363218 210086 363454
rect 209850 362898 210086 363134
rect 240570 363218 240806 363454
rect 240570 362898 240806 363134
rect 71610 331718 71846 331954
rect 71610 331398 71846 331634
rect 102330 331718 102566 331954
rect 102330 331398 102566 331634
rect 133050 331718 133286 331954
rect 133050 331398 133286 331634
rect 163770 331718 164006 331954
rect 163770 331398 164006 331634
rect 194490 331718 194726 331954
rect 194490 331398 194726 331634
rect 225210 331718 225446 331954
rect 225210 331398 225446 331634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 56250 327218 56486 327454
rect 56250 326898 56486 327134
rect 86970 327218 87206 327454
rect 86970 326898 87206 327134
rect 117690 327218 117926 327454
rect 117690 326898 117926 327134
rect 148410 327218 148646 327454
rect 148410 326898 148646 327134
rect 179130 327218 179366 327454
rect 179130 326898 179366 327134
rect 209850 327218 210086 327454
rect 209850 326898 210086 327134
rect 240570 327218 240806 327454
rect 240570 326898 240806 327134
rect 71610 295718 71846 295954
rect 71610 295398 71846 295634
rect 102330 295718 102566 295954
rect 102330 295398 102566 295634
rect 133050 295718 133286 295954
rect 133050 295398 133286 295634
rect 163770 295718 164006 295954
rect 163770 295398 164006 295634
rect 194490 295718 194726 295954
rect 194490 295398 194726 295634
rect 225210 295718 225446 295954
rect 225210 295398 225446 295634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 56250 291218 56486 291454
rect 56250 290898 56486 291134
rect 86970 291218 87206 291454
rect 86970 290898 87206 291134
rect 117690 291218 117926 291454
rect 117690 290898 117926 291134
rect 148410 291218 148646 291454
rect 148410 290898 148646 291134
rect 179130 291218 179366 291454
rect 179130 290898 179366 291134
rect 209850 291218 210086 291454
rect 209850 290898 210086 291134
rect 240570 291218 240806 291454
rect 240570 290898 240806 291134
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 79610 187718 79846 187954
rect 79610 187398 79846 187634
rect 110330 187718 110566 187954
rect 110330 187398 110566 187634
rect 141050 187718 141286 187954
rect 141050 187398 141286 187634
rect 171770 187718 172006 187954
rect 171770 187398 172006 187634
rect 202490 187718 202726 187954
rect 202490 187398 202726 187634
rect 64250 183218 64486 183454
rect 64250 182898 64486 183134
rect 94970 183218 95206 183454
rect 94970 182898 95206 183134
rect 125690 183218 125926 183454
rect 125690 182898 125926 183134
rect 156410 183218 156646 183454
rect 156410 182898 156646 183134
rect 187130 183218 187366 183454
rect 187130 182898 187366 183134
rect 217850 183218 218086 183454
rect 217850 182898 218086 183134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 79610 151718 79846 151954
rect 79610 151398 79846 151634
rect 110330 151718 110566 151954
rect 110330 151398 110566 151634
rect 141050 151718 141286 151954
rect 141050 151398 141286 151634
rect 171770 151718 172006 151954
rect 171770 151398 172006 151634
rect 202490 151718 202726 151954
rect 202490 151398 202726 151634
rect 64250 147218 64486 147454
rect 64250 146898 64486 147134
rect 94970 147218 95206 147454
rect 94970 146898 95206 147134
rect 125690 147218 125926 147454
rect 125690 146898 125926 147134
rect 156410 147218 156646 147454
rect 156410 146898 156646 147134
rect 187130 147218 187366 147454
rect 187130 146898 187366 147134
rect 217850 147218 218086 147454
rect 217850 146898 218086 147134
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 79610 115718 79846 115954
rect 79610 115398 79846 115634
rect 110330 115718 110566 115954
rect 110330 115398 110566 115634
rect 141050 115718 141286 115954
rect 141050 115398 141286 115634
rect 171770 115718 172006 115954
rect 171770 115398 172006 115634
rect 202490 115718 202726 115954
rect 202490 115398 202726 115634
rect 64250 111218 64486 111454
rect 64250 110898 64486 111134
rect 94970 111218 95206 111454
rect 94970 110898 95206 111134
rect 125690 111218 125926 111454
rect 125690 110898 125926 111134
rect 156410 111218 156646 111454
rect 156410 110898 156646 111134
rect 187130 111218 187366 111454
rect 187130 110898 187366 111134
rect 217850 111218 218086 111454
rect 217850 110898 218086 111134
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 79610 79718 79846 79954
rect 79610 79398 79846 79634
rect 110330 79718 110566 79954
rect 110330 79398 110566 79634
rect 141050 79718 141286 79954
rect 141050 79398 141286 79634
rect 171770 79718 172006 79954
rect 171770 79398 172006 79634
rect 202490 79718 202726 79954
rect 202490 79398 202726 79634
rect 64250 75218 64486 75454
rect 64250 74898 64486 75134
rect 94970 75218 95206 75454
rect 94970 74898 95206 75134
rect 125690 75218 125926 75454
rect 125690 74898 125926 75134
rect 156410 75218 156646 75454
rect 156410 74898 156646 75134
rect 187130 75218 187366 75454
rect 187130 74898 187366 75134
rect 217850 75218 218086 75454
rect 217850 74898 218086 75134
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 280826 642125 281062 642361
rect 281146 642125 281382 642361
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 284250 615218 284486 615454
rect 284250 614898 284486 615134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 299610 619718 299846 619954
rect 299610 619398 299846 619634
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 284250 507218 284486 507454
rect 284250 506898 284486 507134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 299610 511718 299846 511954
rect 299610 511398 299846 511634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 316826 642125 317062 642361
rect 317146 642125 317382 642361
rect 314970 615218 315206 615454
rect 314970 614898 315206 615134
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 314970 507218 315206 507454
rect 314970 506898 315206 507134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 304250 327003 304486 327239
rect 334970 327003 335206 327239
rect 319610 295718 319846 295954
rect 319610 295398 319846 295634
rect 304250 291218 304486 291454
rect 304250 290898 304486 291134
rect 334970 291218 335206 291454
rect 334970 290898 335206 291134
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 319610 187718 319846 187954
rect 319610 187398 319846 187634
rect 304250 183218 304486 183454
rect 304250 182898 304486 183134
rect 334970 183218 335206 183454
rect 334970 182898 335206 183134
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 319610 151718 319846 151954
rect 319610 151398 319846 151634
rect 304250 147218 304486 147454
rect 304250 146898 304486 147134
rect 334970 147218 335206 147454
rect 334970 146898 335206 147134
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 319610 115718 319846 115954
rect 319610 115398 319846 115634
rect 304250 111218 304486 111454
rect 304250 110898 304486 111134
rect 334970 111218 335206 111454
rect 334970 110898 335206 111134
rect 319610 79718 319846 79954
rect 319610 79398 319846 79634
rect 304250 75218 304486 75454
rect 304250 74898 304486 75134
rect 334970 75218 335206 75454
rect 334970 74898 335206 75134
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642125 389062 642361
rect 389146 642125 389382 642361
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 379610 619718 379846 619954
rect 379610 619398 379846 619634
rect 364250 615218 364486 615454
rect 364250 614898 364486 615134
rect 394970 615218 395206 615454
rect 394970 614898 395206 615134
rect 364250 543218 364486 543454
rect 364250 542898 364486 543134
rect 364250 507218 364486 507454
rect 364250 506898 364486 507134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552125 371062 552361
rect 371146 552125 371382 552361
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379610 511718 379846 511954
rect 379610 511398 379846 511634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 394970 543218 395206 543454
rect 394970 542898 395206 543134
rect 394970 507218 395206 507454
rect 394970 506898 395206 507134
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 484250 615218 484486 615454
rect 484250 614898 484486 615134
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 487934 511718 488170 511954
rect 487934 511398 488170 511634
rect 484460 507218 484696 507454
rect 484460 506898 484696 507134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 494882 511718 495118 511954
rect 494882 511398 495118 511634
rect 491408 507218 491644 507454
rect 491408 506898 491644 507134
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 496826 642125 497062 642361
rect 497146 642125 497382 642361
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 499610 619718 499846 619954
rect 499610 619398 499846 619634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 501830 511718 502066 511954
rect 501830 511398 502066 511634
rect 498356 507218 498592 507454
rect 498356 506898 498592 507134
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 505304 507218 505540 507454
rect 505304 506898 505540 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 514970 615218 515206 615454
rect 514970 614898 515206 615134
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 71610 655954
rect 71846 655718 102330 655954
rect 102566 655718 133050 655954
rect 133286 655718 163770 655954
rect 164006 655718 194490 655954
rect 194726 655718 225210 655954
rect 225446 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 71610 655634
rect 71846 655398 102330 655634
rect 102566 655398 133050 655634
rect 133286 655398 163770 655634
rect 164006 655398 194490 655634
rect 194726 655398 225210 655634
rect 225446 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 56250 651454
rect 56486 651218 86970 651454
rect 87206 651218 117690 651454
rect 117926 651218 148410 651454
rect 148646 651218 179130 651454
rect 179366 651218 209850 651454
rect 210086 651218 240570 651454
rect 240806 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 56250 651134
rect 56486 650898 86970 651134
rect 87206 650898 117690 651134
rect 117926 650898 148410 651134
rect 148646 650898 179130 651134
rect 179366 650898 209850 651134
rect 210086 650898 240570 651134
rect 240806 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642361 352826 642454
rect 29382 642218 280826 642361
rect -8726 642134 280826 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 642125 280826 642134
rect 281062 642125 281146 642361
rect 281382 642125 316826 642361
rect 317062 642125 317146 642361
rect 317382 642218 352826 642361
rect 353062 642218 353146 642454
rect 353382 642361 424826 642454
rect 353382 642218 388826 642361
rect 317382 642134 388826 642218
rect 317382 642125 352826 642134
rect 29382 641898 352826 642125
rect 353062 641898 353146 642134
rect 353382 642125 388826 642134
rect 389062 642125 389146 642361
rect 389382 642218 424826 642361
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642361 532826 642454
rect 461382 642218 496826 642361
rect 389382 642134 496826 642218
rect 389382 642125 424826 642134
rect 353382 641898 424826 642125
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 642125 496826 642134
rect 497062 642125 497146 642361
rect 497382 642218 532826 642361
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect 497382 642134 592650 642218
rect 497382 642125 532826 642134
rect 461382 641898 532826 642125
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 71610 619954
rect 71846 619718 102330 619954
rect 102566 619718 133050 619954
rect 133286 619718 163770 619954
rect 164006 619718 194490 619954
rect 194726 619718 225210 619954
rect 225446 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 299610 619954
rect 299846 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 379610 619954
rect 379846 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 499610 619954
rect 499846 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 71610 619634
rect 71846 619398 102330 619634
rect 102566 619398 133050 619634
rect 133286 619398 163770 619634
rect 164006 619398 194490 619634
rect 194726 619398 225210 619634
rect 225446 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 299610 619634
rect 299846 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 379610 619634
rect 379846 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 499610 619634
rect 499846 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 56250 615454
rect 56486 615218 86970 615454
rect 87206 615218 117690 615454
rect 117926 615218 148410 615454
rect 148646 615218 179130 615454
rect 179366 615218 209850 615454
rect 210086 615218 240570 615454
rect 240806 615218 284250 615454
rect 284486 615218 314970 615454
rect 315206 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 364250 615454
rect 364486 615218 394970 615454
rect 395206 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 484250 615454
rect 484486 615218 514970 615454
rect 515206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 56250 615134
rect 56486 614898 86970 615134
rect 87206 614898 117690 615134
rect 117926 614898 148410 615134
rect 148646 614898 179130 615134
rect 179366 614898 209850 615134
rect 210086 614898 240570 615134
rect 240806 614898 284250 615134
rect 284486 614898 314970 615134
rect 315206 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 364250 615134
rect 364486 614898 394970 615134
rect 395206 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 484250 615134
rect 484486 614898 514970 615134
rect 515206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 71610 583954
rect 71846 583718 102330 583954
rect 102566 583718 133050 583954
rect 133286 583718 163770 583954
rect 164006 583718 194490 583954
rect 194726 583718 225210 583954
rect 225446 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 71610 583634
rect 71846 583398 102330 583634
rect 102566 583398 133050 583634
rect 133286 583398 163770 583634
rect 164006 583398 194490 583634
rect 194726 583398 225210 583634
rect 225446 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 56250 579454
rect 56486 579218 86970 579454
rect 87206 579218 117690 579454
rect 117926 579218 148410 579454
rect 148646 579218 179130 579454
rect 179366 579218 209850 579454
rect 210086 579218 240570 579454
rect 240806 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 56250 579134
rect 56486 578898 86970 579134
rect 87206 578898 117690 579134
rect 117926 578898 148410 579134
rect 148646 578898 179130 579134
rect 179366 578898 209850 579134
rect 210086 578898 240570 579134
rect 240806 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552361 406826 552454
rect 335382 552218 370826 552361
rect -8726 552134 370826 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 552125 370826 552134
rect 371062 552125 371146 552361
rect 371382 552218 406826 552361
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect 371382 552134 592650 552218
rect 371382 552125 406826 552134
rect 335382 551898 406826 552125
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 71610 547954
rect 71846 547718 102330 547954
rect 102566 547718 133050 547954
rect 133286 547718 163770 547954
rect 164006 547718 194490 547954
rect 194726 547718 225210 547954
rect 225446 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 71610 547634
rect 71846 547398 102330 547634
rect 102566 547398 133050 547634
rect 133286 547398 163770 547634
rect 164006 547398 194490 547634
rect 194726 547398 225210 547634
rect 225446 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 56250 543454
rect 56486 543218 86970 543454
rect 87206 543218 117690 543454
rect 117926 543218 148410 543454
rect 148646 543218 179130 543454
rect 179366 543218 209850 543454
rect 210086 543218 240570 543454
rect 240806 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 364250 543454
rect 364486 543218 394970 543454
rect 395206 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 56250 543134
rect 56486 542898 86970 543134
rect 87206 542898 117690 543134
rect 117926 542898 148410 543134
rect 148646 542898 179130 543134
rect 179366 542898 209850 543134
rect 210086 542898 240570 543134
rect 240806 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 364250 543134
rect 364486 542898 394970 543134
rect 395206 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 71610 511954
rect 71846 511718 102330 511954
rect 102566 511718 133050 511954
rect 133286 511718 163770 511954
rect 164006 511718 194490 511954
rect 194726 511718 225210 511954
rect 225446 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 299610 511954
rect 299846 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 379610 511954
rect 379846 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 487934 511954
rect 488170 511718 494882 511954
rect 495118 511718 501830 511954
rect 502066 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 71610 511634
rect 71846 511398 102330 511634
rect 102566 511398 133050 511634
rect 133286 511398 163770 511634
rect 164006 511398 194490 511634
rect 194726 511398 225210 511634
rect 225446 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 299610 511634
rect 299846 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 379610 511634
rect 379846 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 487934 511634
rect 488170 511398 494882 511634
rect 495118 511398 501830 511634
rect 502066 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 56250 507454
rect 56486 507218 86970 507454
rect 87206 507218 117690 507454
rect 117926 507218 148410 507454
rect 148646 507218 179130 507454
rect 179366 507218 209850 507454
rect 210086 507218 240570 507454
rect 240806 507218 284250 507454
rect 284486 507218 314970 507454
rect 315206 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 364250 507454
rect 364486 507218 394970 507454
rect 395206 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 484460 507454
rect 484696 507218 491408 507454
rect 491644 507218 498356 507454
rect 498592 507218 505304 507454
rect 505540 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 56250 507134
rect 56486 506898 86970 507134
rect 87206 506898 117690 507134
rect 117926 506898 148410 507134
rect 148646 506898 179130 507134
rect 179366 506898 209850 507134
rect 210086 506898 240570 507134
rect 240806 506898 284250 507134
rect 284486 506898 314970 507134
rect 315206 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 364250 507134
rect 364486 506898 394970 507134
rect 395206 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 484460 507134
rect 484696 506898 491408 507134
rect 491644 506898 498356 507134
rect 498592 506898 505304 507134
rect 505540 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 71610 475954
rect 71846 475718 102330 475954
rect 102566 475718 133050 475954
rect 133286 475718 163770 475954
rect 164006 475718 194490 475954
rect 194726 475718 225210 475954
rect 225446 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 71610 475634
rect 71846 475398 102330 475634
rect 102566 475398 133050 475634
rect 133286 475398 163770 475634
rect 164006 475398 194490 475634
rect 194726 475398 225210 475634
rect 225446 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 56250 471454
rect 56486 471218 86970 471454
rect 87206 471218 117690 471454
rect 117926 471218 148410 471454
rect 148646 471218 179130 471454
rect 179366 471218 209850 471454
rect 210086 471218 240570 471454
rect 240806 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 56250 471134
rect 56486 470898 86970 471134
rect 87206 470898 117690 471134
rect 117926 470898 148410 471134
rect 148646 470898 179130 471134
rect 179366 470898 209850 471134
rect 210086 470898 240570 471134
rect 240806 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 71610 439954
rect 71846 439718 102330 439954
rect 102566 439718 133050 439954
rect 133286 439718 163770 439954
rect 164006 439718 194490 439954
rect 194726 439718 225210 439954
rect 225446 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 71610 439634
rect 71846 439398 102330 439634
rect 102566 439398 133050 439634
rect 133286 439398 163770 439634
rect 164006 439398 194490 439634
rect 194726 439398 225210 439634
rect 225446 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 56250 435454
rect 56486 435218 86970 435454
rect 87206 435218 117690 435454
rect 117926 435218 148410 435454
rect 148646 435218 179130 435454
rect 179366 435218 209850 435454
rect 210086 435218 240570 435454
rect 240806 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 56250 435134
rect 56486 434898 86970 435134
rect 87206 434898 117690 435134
rect 117926 434898 148410 435134
rect 148646 434898 179130 435134
rect 179366 434898 209850 435134
rect 210086 434898 240570 435134
rect 240806 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 71610 403954
rect 71846 403718 102330 403954
rect 102566 403718 133050 403954
rect 133286 403718 163770 403954
rect 164006 403718 194490 403954
rect 194726 403718 225210 403954
rect 225446 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 71610 403634
rect 71846 403398 102330 403634
rect 102566 403398 133050 403634
rect 133286 403398 163770 403634
rect 164006 403398 194490 403634
rect 194726 403398 225210 403634
rect 225446 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 56250 399454
rect 56486 399218 86970 399454
rect 87206 399218 117690 399454
rect 117926 399218 148410 399454
rect 148646 399218 179130 399454
rect 179366 399218 209850 399454
rect 210086 399218 240570 399454
rect 240806 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 56250 399134
rect 56486 398898 86970 399134
rect 87206 398898 117690 399134
rect 117926 398898 148410 399134
rect 148646 398898 179130 399134
rect 179366 398898 209850 399134
rect 210086 398898 240570 399134
rect 240806 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 71610 367954
rect 71846 367718 102330 367954
rect 102566 367718 133050 367954
rect 133286 367718 163770 367954
rect 164006 367718 194490 367954
rect 194726 367718 225210 367954
rect 225446 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 71610 367634
rect 71846 367398 102330 367634
rect 102566 367398 133050 367634
rect 133286 367398 163770 367634
rect 164006 367398 194490 367634
rect 194726 367398 225210 367634
rect 225446 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 56250 363454
rect 56486 363218 86970 363454
rect 87206 363218 117690 363454
rect 117926 363218 148410 363454
rect 148646 363218 179130 363454
rect 179366 363218 209850 363454
rect 210086 363218 240570 363454
rect 240806 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 56250 363134
rect 56486 362898 86970 363134
rect 87206 362898 117690 363134
rect 117926 362898 148410 363134
rect 148646 362898 179130 363134
rect 179366 362898 209850 363134
rect 210086 362898 240570 363134
rect 240806 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 71610 331954
rect 71846 331718 102330 331954
rect 102566 331718 133050 331954
rect 133286 331718 163770 331954
rect 164006 331718 194490 331954
rect 194726 331718 225210 331954
rect 225446 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 71610 331634
rect 71846 331398 102330 331634
rect 102566 331398 133050 331634
rect 133286 331398 163770 331634
rect 164006 331398 194490 331634
rect 194726 331398 225210 331634
rect 225446 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 56250 327454
rect 56486 327218 86970 327454
rect 87206 327218 117690 327454
rect 117926 327218 148410 327454
rect 148646 327218 179130 327454
rect 179366 327218 209850 327454
rect 210086 327218 240570 327454
rect 240806 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327239 361826 327454
rect 290382 327218 304250 327239
rect -8726 327134 304250 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 56250 327134
rect 56486 326898 86970 327134
rect 87206 326898 117690 327134
rect 117926 326898 148410 327134
rect 148646 326898 179130 327134
rect 179366 326898 209850 327134
rect 210086 326898 240570 327134
rect 240806 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 327003 304250 327134
rect 304486 327003 334970 327239
rect 335206 327218 361826 327239
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect 335206 327134 592650 327218
rect 335206 327003 361826 327134
rect 290382 326898 361826 327003
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 71610 295954
rect 71846 295718 102330 295954
rect 102566 295718 133050 295954
rect 133286 295718 163770 295954
rect 164006 295718 194490 295954
rect 194726 295718 225210 295954
rect 225446 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 319610 295954
rect 319846 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 71610 295634
rect 71846 295398 102330 295634
rect 102566 295398 133050 295634
rect 133286 295398 163770 295634
rect 164006 295398 194490 295634
rect 194726 295398 225210 295634
rect 225446 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 319610 295634
rect 319846 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 56250 291454
rect 56486 291218 86970 291454
rect 87206 291218 117690 291454
rect 117926 291218 148410 291454
rect 148646 291218 179130 291454
rect 179366 291218 209850 291454
rect 210086 291218 240570 291454
rect 240806 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 304250 291454
rect 304486 291218 334970 291454
rect 335206 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 56250 291134
rect 56486 290898 86970 291134
rect 87206 290898 117690 291134
rect 117926 290898 148410 291134
rect 148646 290898 179130 291134
rect 179366 290898 209850 291134
rect 210086 290898 240570 291134
rect 240806 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 304250 291134
rect 304486 290898 334970 291134
rect 335206 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 79610 187954
rect 79846 187718 110330 187954
rect 110566 187718 141050 187954
rect 141286 187718 171770 187954
rect 172006 187718 202490 187954
rect 202726 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 319610 187954
rect 319846 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 79610 187634
rect 79846 187398 110330 187634
rect 110566 187398 141050 187634
rect 141286 187398 171770 187634
rect 172006 187398 202490 187634
rect 202726 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 319610 187634
rect 319846 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 64250 183454
rect 64486 183218 94970 183454
rect 95206 183218 125690 183454
rect 125926 183218 156410 183454
rect 156646 183218 187130 183454
rect 187366 183218 217850 183454
rect 218086 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 304250 183454
rect 304486 183218 334970 183454
rect 335206 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 64250 183134
rect 64486 182898 94970 183134
rect 95206 182898 125690 183134
rect 125926 182898 156410 183134
rect 156646 182898 187130 183134
rect 187366 182898 217850 183134
rect 218086 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 304250 183134
rect 304486 182898 334970 183134
rect 335206 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 79610 151954
rect 79846 151718 110330 151954
rect 110566 151718 141050 151954
rect 141286 151718 171770 151954
rect 172006 151718 202490 151954
rect 202726 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 319610 151954
rect 319846 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 79610 151634
rect 79846 151398 110330 151634
rect 110566 151398 141050 151634
rect 141286 151398 171770 151634
rect 172006 151398 202490 151634
rect 202726 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 319610 151634
rect 319846 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 64250 147454
rect 64486 147218 94970 147454
rect 95206 147218 125690 147454
rect 125926 147218 156410 147454
rect 156646 147218 187130 147454
rect 187366 147218 217850 147454
rect 218086 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 304250 147454
rect 304486 147218 334970 147454
rect 335206 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 64250 147134
rect 64486 146898 94970 147134
rect 95206 146898 125690 147134
rect 125926 146898 156410 147134
rect 156646 146898 187130 147134
rect 187366 146898 217850 147134
rect 218086 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 304250 147134
rect 304486 146898 334970 147134
rect 335206 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 79610 115954
rect 79846 115718 110330 115954
rect 110566 115718 141050 115954
rect 141286 115718 171770 115954
rect 172006 115718 202490 115954
rect 202726 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 319610 115954
rect 319846 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 79610 115634
rect 79846 115398 110330 115634
rect 110566 115398 141050 115634
rect 141286 115398 171770 115634
rect 172006 115398 202490 115634
rect 202726 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 319610 115634
rect 319846 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 64250 111454
rect 64486 111218 94970 111454
rect 95206 111218 125690 111454
rect 125926 111218 156410 111454
rect 156646 111218 187130 111454
rect 187366 111218 217850 111454
rect 218086 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 304250 111454
rect 304486 111218 334970 111454
rect 335206 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 64250 111134
rect 64486 110898 94970 111134
rect 95206 110898 125690 111134
rect 125926 110898 156410 111134
rect 156646 110898 187130 111134
rect 187366 110898 217850 111134
rect 218086 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 304250 111134
rect 304486 110898 334970 111134
rect 335206 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 79610 79954
rect 79846 79718 110330 79954
rect 110566 79718 141050 79954
rect 141286 79718 171770 79954
rect 172006 79718 202490 79954
rect 202726 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 319610 79954
rect 319846 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 79610 79634
rect 79846 79398 110330 79634
rect 110566 79398 141050 79634
rect 141286 79398 171770 79634
rect 172006 79398 202490 79634
rect 202726 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 319610 79634
rect 319846 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 64250 75454
rect 64486 75218 94970 75454
rect 95206 75218 125690 75454
rect 125926 75218 156410 75454
rect 156646 75218 187130 75454
rect 187366 75218 217850 75454
rect 218086 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 304250 75454
rect 304486 75218 334970 75454
rect 335206 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 64250 75134
rect 64486 74898 94970 75134
rect 95206 74898 125690 75134
rect 125926 74898 156410 75134
rect 156646 74898 187130 75134
rect 187366 74898 217850 75134
rect 218086 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 304250 75134
rect 304486 74898 334970 75134
rect 335206 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use clock_div  top_cw.clock_div
timestamp 0
transform 1 0 480000 0 1 600000
box 0 0 40000 40000
use top_cw_logic  top_cw.top_cw_logic
timestamp 0
transform 1 0 360000 0 1 500000
box 0 0 40000 50000
use core  top_cw.upc.core
timestamp 0
transform 1 0 300000 0 1 60000
box 0 2048 40000 160000
use dcache  top_cw.upc.dcache
timestamp 0
transform 1 0 52000 0 1 280000
box 0 2128 200000 379760
use icache  top_cw.upc.icache
timestamp 0
transform 1 0 60000 0 1 60000
box 0 2042 160000 157808
use upper_core_logic  top_cw.upc.upper_core_logic
timestamp 0
transform 1 0 300000 0 1 280000
box 0 0 50000 50000
use wishbone_arbiter  top_cw.upc.wb_arbiter
timestamp 0
transform 1 0 280000 0 1 500000
box 1066 0 40000 40000
use wb_compressor  top_cw.wb_compressor
timestamp 0
transform 1 0 280000 0 1 600000
box 0 0 39362 40000
use wb_cross_clk  top_cw.wb_cross_clk
timestamp 0
transform 1 0 360000 0 1 600000
box 1066 0 38862 40000
use uprj_w_const  uprj_w_const
timestamp 0
transform 1 0 480000 0 1 500000
box 0 0 30000 30000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 664000 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 664000 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 664000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 664000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 664000 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 278000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 664000 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 542000 290414 598000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 642000 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 332000 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 642000 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 642000 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 532000 506414 598000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 642000 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 222000 83414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 664000 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 222000 119414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 664000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 222000 155414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 664000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 222000 191414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 664000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 664000 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 222000 299414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 332000 299414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 542000 299414 598000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 642000 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 222000 335414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 332000 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 552000 371414 598000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 642000 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 532000 479414 598000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 642000 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 598000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 642000 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 222000 56414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 664000 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 222000 92414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 664000 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 222000 128414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 664000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 222000 164414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 664000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 222000 200414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 664000 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 664000 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 222000 308414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 332000 308414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 542000 308414 598000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 642000 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 222000 344414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 332000 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 552000 380414 598000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 642000 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 532000 488414 598000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 642000 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 598000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 642000 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 664000 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 664000 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 664000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 664000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 664000 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 278000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 664000 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 642000 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 332000 317414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 642000 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 278000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 332000 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 642000 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 532000 497414 598000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 642000 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 222000 60914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 664000 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 222000 96914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 664000 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 222000 132914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 664000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 222000 168914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 664000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 222000 204914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 664000 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 664000 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 642000 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 222000 312914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 332000 312914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 642000 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 332000 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 642000 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 642000 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 664000 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 664000 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 664000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 664000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 664000 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 278000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 664000 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 642000 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 332000 321914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 642000 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 642000 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 642000 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 532000 501914 598000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 642000 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 222000 78914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 664000 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 222000 114914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 664000 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 222000 150914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 664000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 222000 186914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 664000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 222000 222914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 664000 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 542000 294914 598000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 642000 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 222000 330914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 332000 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 642000 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 642000 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 532000 510914 598000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 642000 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 664000 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 222000 87914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 664000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 222000 123914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 664000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 222000 159914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 664000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 222000 195914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 664000 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 664000 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 222000 303914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 332000 303914 498000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 542000 303914 598000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 642000 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 222000 339914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 332000 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 498000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 552000 375914 598000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 642000 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 498000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 532000 483914 598000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 642000 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 598000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 642000 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
