VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO interconnect_inner
  CLASS BLOCK ;
  FOREIGN interconnect_inner ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 800.000 ;
  PIN c0_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END c0_clk
  PIN c0_dbg_pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END c0_dbg_pc[0]
  PIN c0_dbg_pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END c0_dbg_pc[10]
  PIN c0_dbg_pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END c0_dbg_pc[11]
  PIN c0_dbg_pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END c0_dbg_pc[12]
  PIN c0_dbg_pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END c0_dbg_pc[13]
  PIN c0_dbg_pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END c0_dbg_pc[14]
  PIN c0_dbg_pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END c0_dbg_pc[15]
  PIN c0_dbg_pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END c0_dbg_pc[1]
  PIN c0_dbg_pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END c0_dbg_pc[2]
  PIN c0_dbg_pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END c0_dbg_pc[3]
  PIN c0_dbg_pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END c0_dbg_pc[4]
  PIN c0_dbg_pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END c0_dbg_pc[5]
  PIN c0_dbg_pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END c0_dbg_pc[6]
  PIN c0_dbg_pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END c0_dbg_pc[7]
  PIN c0_dbg_pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END c0_dbg_pc[8]
  PIN c0_dbg_pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END c0_dbg_pc[9]
  PIN c0_dbg_r0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END c0_dbg_r0[0]
  PIN c0_dbg_r0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END c0_dbg_r0[10]
  PIN c0_dbg_r0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END c0_dbg_r0[11]
  PIN c0_dbg_r0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END c0_dbg_r0[12]
  PIN c0_dbg_r0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END c0_dbg_r0[13]
  PIN c0_dbg_r0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END c0_dbg_r0[14]
  PIN c0_dbg_r0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END c0_dbg_r0[15]
  PIN c0_dbg_r0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END c0_dbg_r0[1]
  PIN c0_dbg_r0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END c0_dbg_r0[2]
  PIN c0_dbg_r0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END c0_dbg_r0[3]
  PIN c0_dbg_r0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END c0_dbg_r0[4]
  PIN c0_dbg_r0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END c0_dbg_r0[5]
  PIN c0_dbg_r0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END c0_dbg_r0[6]
  PIN c0_dbg_r0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END c0_dbg_r0[7]
  PIN c0_dbg_r0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END c0_dbg_r0[8]
  PIN c0_dbg_r0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END c0_dbg_r0[9]
  PIN c0_disable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END c0_disable
  PIN c0_i_core_int_sreg[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END c0_i_core_int_sreg[0]
  PIN c0_i_core_int_sreg[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END c0_i_core_int_sreg[10]
  PIN c0_i_core_int_sreg[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END c0_i_core_int_sreg[11]
  PIN c0_i_core_int_sreg[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END c0_i_core_int_sreg[12]
  PIN c0_i_core_int_sreg[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END c0_i_core_int_sreg[13]
  PIN c0_i_core_int_sreg[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END c0_i_core_int_sreg[14]
  PIN c0_i_core_int_sreg[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END c0_i_core_int_sreg[15]
  PIN c0_i_core_int_sreg[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END c0_i_core_int_sreg[1]
  PIN c0_i_core_int_sreg[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END c0_i_core_int_sreg[2]
  PIN c0_i_core_int_sreg[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END c0_i_core_int_sreg[3]
  PIN c0_i_core_int_sreg[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END c0_i_core_int_sreg[4]
  PIN c0_i_core_int_sreg[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END c0_i_core_int_sreg[5]
  PIN c0_i_core_int_sreg[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END c0_i_core_int_sreg[6]
  PIN c0_i_core_int_sreg[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END c0_i_core_int_sreg[7]
  PIN c0_i_core_int_sreg[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END c0_i_core_int_sreg[8]
  PIN c0_i_core_int_sreg[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END c0_i_core_int_sreg[9]
  PIN c0_i_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END c0_i_irq
  PIN c0_i_mc_core_int
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END c0_i_mc_core_int
  PIN c0_i_mem_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END c0_i_mem_ack
  PIN c0_i_mem_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END c0_i_mem_data[0]
  PIN c0_i_mem_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END c0_i_mem_data[10]
  PIN c0_i_mem_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END c0_i_mem_data[11]
  PIN c0_i_mem_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END c0_i_mem_data[12]
  PIN c0_i_mem_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END c0_i_mem_data[13]
  PIN c0_i_mem_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END c0_i_mem_data[14]
  PIN c0_i_mem_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END c0_i_mem_data[15]
  PIN c0_i_mem_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END c0_i_mem_data[1]
  PIN c0_i_mem_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END c0_i_mem_data[2]
  PIN c0_i_mem_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END c0_i_mem_data[3]
  PIN c0_i_mem_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END c0_i_mem_data[4]
  PIN c0_i_mem_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END c0_i_mem_data[5]
  PIN c0_i_mem_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END c0_i_mem_data[6]
  PIN c0_i_mem_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END c0_i_mem_data[7]
  PIN c0_i_mem_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END c0_i_mem_data[8]
  PIN c0_i_mem_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END c0_i_mem_data[9]
  PIN c0_i_mem_exception
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END c0_i_mem_exception
  PIN c0_i_req_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END c0_i_req_data[0]
  PIN c0_i_req_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END c0_i_req_data[10]
  PIN c0_i_req_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END c0_i_req_data[11]
  PIN c0_i_req_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END c0_i_req_data[12]
  PIN c0_i_req_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END c0_i_req_data[13]
  PIN c0_i_req_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END c0_i_req_data[14]
  PIN c0_i_req_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END c0_i_req_data[15]
  PIN c0_i_req_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END c0_i_req_data[16]
  PIN c0_i_req_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END c0_i_req_data[17]
  PIN c0_i_req_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END c0_i_req_data[18]
  PIN c0_i_req_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END c0_i_req_data[19]
  PIN c0_i_req_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END c0_i_req_data[1]
  PIN c0_i_req_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END c0_i_req_data[20]
  PIN c0_i_req_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END c0_i_req_data[21]
  PIN c0_i_req_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END c0_i_req_data[22]
  PIN c0_i_req_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END c0_i_req_data[23]
  PIN c0_i_req_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END c0_i_req_data[24]
  PIN c0_i_req_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END c0_i_req_data[25]
  PIN c0_i_req_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END c0_i_req_data[26]
  PIN c0_i_req_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END c0_i_req_data[27]
  PIN c0_i_req_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END c0_i_req_data[28]
  PIN c0_i_req_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END c0_i_req_data[29]
  PIN c0_i_req_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END c0_i_req_data[2]
  PIN c0_i_req_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END c0_i_req_data[30]
  PIN c0_i_req_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END c0_i_req_data[31]
  PIN c0_i_req_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END c0_i_req_data[3]
  PIN c0_i_req_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END c0_i_req_data[4]
  PIN c0_i_req_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END c0_i_req_data[5]
  PIN c0_i_req_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END c0_i_req_data[6]
  PIN c0_i_req_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END c0_i_req_data[7]
  PIN c0_i_req_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END c0_i_req_data[8]
  PIN c0_i_req_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END c0_i_req_data[9]
  PIN c0_i_req_data_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END c0_i_req_data_valid
  PIN c0_o_c_data_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END c0_o_c_data_page
  PIN c0_o_c_instr_long
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END c0_o_c_instr_long
  PIN c0_o_c_instr_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END c0_o_c_instr_page
  PIN c0_o_icache_flush
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END c0_o_icache_flush
  PIN c0_o_instr_long_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END c0_o_instr_long_addr[0]
  PIN c0_o_instr_long_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END c0_o_instr_long_addr[1]
  PIN c0_o_instr_long_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END c0_o_instr_long_addr[2]
  PIN c0_o_instr_long_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END c0_o_instr_long_addr[3]
  PIN c0_o_instr_long_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END c0_o_instr_long_addr[4]
  PIN c0_o_instr_long_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END c0_o_instr_long_addr[5]
  PIN c0_o_instr_long_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END c0_o_instr_long_addr[6]
  PIN c0_o_instr_long_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END c0_o_instr_long_addr[7]
  PIN c0_o_mem_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END c0_o_mem_addr[0]
  PIN c0_o_mem_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END c0_o_mem_addr[10]
  PIN c0_o_mem_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END c0_o_mem_addr[11]
  PIN c0_o_mem_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END c0_o_mem_addr[12]
  PIN c0_o_mem_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END c0_o_mem_addr[13]
  PIN c0_o_mem_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END c0_o_mem_addr[14]
  PIN c0_o_mem_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END c0_o_mem_addr[15]
  PIN c0_o_mem_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END c0_o_mem_addr[1]
  PIN c0_o_mem_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END c0_o_mem_addr[2]
  PIN c0_o_mem_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END c0_o_mem_addr[3]
  PIN c0_o_mem_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END c0_o_mem_addr[4]
  PIN c0_o_mem_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END c0_o_mem_addr[5]
  PIN c0_o_mem_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END c0_o_mem_addr[6]
  PIN c0_o_mem_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END c0_o_mem_addr[7]
  PIN c0_o_mem_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END c0_o_mem_addr[8]
  PIN c0_o_mem_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END c0_o_mem_addr[9]
  PIN c0_o_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END c0_o_mem_data[0]
  PIN c0_o_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END c0_o_mem_data[10]
  PIN c0_o_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END c0_o_mem_data[11]
  PIN c0_o_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END c0_o_mem_data[12]
  PIN c0_o_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END c0_o_mem_data[13]
  PIN c0_o_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END c0_o_mem_data[14]
  PIN c0_o_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END c0_o_mem_data[15]
  PIN c0_o_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END c0_o_mem_data[1]
  PIN c0_o_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END c0_o_mem_data[2]
  PIN c0_o_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END c0_o_mem_data[3]
  PIN c0_o_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END c0_o_mem_data[4]
  PIN c0_o_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END c0_o_mem_data[5]
  PIN c0_o_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END c0_o_mem_data[6]
  PIN c0_o_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END c0_o_mem_data[7]
  PIN c0_o_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END c0_o_mem_data[8]
  PIN c0_o_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END c0_o_mem_data[9]
  PIN c0_o_mem_high_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END c0_o_mem_high_addr[0]
  PIN c0_o_mem_high_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END c0_o_mem_high_addr[1]
  PIN c0_o_mem_high_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END c0_o_mem_high_addr[2]
  PIN c0_o_mem_high_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END c0_o_mem_high_addr[3]
  PIN c0_o_mem_high_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END c0_o_mem_high_addr[4]
  PIN c0_o_mem_high_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END c0_o_mem_high_addr[5]
  PIN c0_o_mem_high_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END c0_o_mem_high_addr[6]
  PIN c0_o_mem_high_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END c0_o_mem_high_addr[7]
  PIN c0_o_mem_long_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END c0_o_mem_long_mode
  PIN c0_o_mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END c0_o_mem_req
  PIN c0_o_mem_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END c0_o_mem_sel[0]
  PIN c0_o_mem_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END c0_o_mem_sel[1]
  PIN c0_o_mem_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END c0_o_mem_we
  PIN c0_o_req_active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END c0_o_req_active
  PIN c0_o_req_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END c0_o_req_addr[0]
  PIN c0_o_req_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END c0_o_req_addr[10]
  PIN c0_o_req_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END c0_o_req_addr[11]
  PIN c0_o_req_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END c0_o_req_addr[12]
  PIN c0_o_req_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END c0_o_req_addr[13]
  PIN c0_o_req_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END c0_o_req_addr[14]
  PIN c0_o_req_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END c0_o_req_addr[15]
  PIN c0_o_req_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END c0_o_req_addr[1]
  PIN c0_o_req_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END c0_o_req_addr[2]
  PIN c0_o_req_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END c0_o_req_addr[3]
  PIN c0_o_req_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END c0_o_req_addr[4]
  PIN c0_o_req_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END c0_o_req_addr[5]
  PIN c0_o_req_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END c0_o_req_addr[6]
  PIN c0_o_req_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END c0_o_req_addr[7]
  PIN c0_o_req_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END c0_o_req_addr[8]
  PIN c0_o_req_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END c0_o_req_addr[9]
  PIN c0_o_req_ppl_submit
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END c0_o_req_ppl_submit
  PIN c0_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END c0_rst
  PIN c0_sr_bus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END c0_sr_bus_addr[0]
  PIN c0_sr_bus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END c0_sr_bus_addr[10]
  PIN c0_sr_bus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END c0_sr_bus_addr[11]
  PIN c0_sr_bus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END c0_sr_bus_addr[12]
  PIN c0_sr_bus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END c0_sr_bus_addr[13]
  PIN c0_sr_bus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END c0_sr_bus_addr[14]
  PIN c0_sr_bus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END c0_sr_bus_addr[15]
  PIN c0_sr_bus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END c0_sr_bus_addr[1]
  PIN c0_sr_bus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END c0_sr_bus_addr[2]
  PIN c0_sr_bus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END c0_sr_bus_addr[3]
  PIN c0_sr_bus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END c0_sr_bus_addr[4]
  PIN c0_sr_bus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END c0_sr_bus_addr[5]
  PIN c0_sr_bus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END c0_sr_bus_addr[6]
  PIN c0_sr_bus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END c0_sr_bus_addr[7]
  PIN c0_sr_bus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END c0_sr_bus_addr[8]
  PIN c0_sr_bus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END c0_sr_bus_addr[9]
  PIN c0_sr_bus_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END c0_sr_bus_data_o[0]
  PIN c0_sr_bus_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END c0_sr_bus_data_o[10]
  PIN c0_sr_bus_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END c0_sr_bus_data_o[11]
  PIN c0_sr_bus_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END c0_sr_bus_data_o[12]
  PIN c0_sr_bus_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END c0_sr_bus_data_o[13]
  PIN c0_sr_bus_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END c0_sr_bus_data_o[14]
  PIN c0_sr_bus_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END c0_sr_bus_data_o[15]
  PIN c0_sr_bus_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END c0_sr_bus_data_o[1]
  PIN c0_sr_bus_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END c0_sr_bus_data_o[2]
  PIN c0_sr_bus_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END c0_sr_bus_data_o[3]
  PIN c0_sr_bus_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END c0_sr_bus_data_o[4]
  PIN c0_sr_bus_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END c0_sr_bus_data_o[5]
  PIN c0_sr_bus_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END c0_sr_bus_data_o[6]
  PIN c0_sr_bus_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END c0_sr_bus_data_o[7]
  PIN c0_sr_bus_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END c0_sr_bus_data_o[8]
  PIN c0_sr_bus_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END c0_sr_bus_data_o[9]
  PIN c0_sr_bus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END c0_sr_bus_we
  PIN c1_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END c1_clk
  PIN c1_dbg_pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END c1_dbg_pc[0]
  PIN c1_dbg_pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END c1_dbg_pc[10]
  PIN c1_dbg_pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END c1_dbg_pc[11]
  PIN c1_dbg_pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END c1_dbg_pc[12]
  PIN c1_dbg_pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END c1_dbg_pc[13]
  PIN c1_dbg_pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END c1_dbg_pc[14]
  PIN c1_dbg_pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END c1_dbg_pc[15]
  PIN c1_dbg_pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END c1_dbg_pc[1]
  PIN c1_dbg_pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END c1_dbg_pc[2]
  PIN c1_dbg_pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END c1_dbg_pc[3]
  PIN c1_dbg_pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END c1_dbg_pc[4]
  PIN c1_dbg_pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END c1_dbg_pc[5]
  PIN c1_dbg_pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END c1_dbg_pc[6]
  PIN c1_dbg_pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END c1_dbg_pc[7]
  PIN c1_dbg_pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END c1_dbg_pc[8]
  PIN c1_dbg_pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END c1_dbg_pc[9]
  PIN c1_dbg_r0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END c1_dbg_r0[0]
  PIN c1_dbg_r0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END c1_dbg_r0[10]
  PIN c1_dbg_r0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END c1_dbg_r0[11]
  PIN c1_dbg_r0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END c1_dbg_r0[12]
  PIN c1_dbg_r0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END c1_dbg_r0[13]
  PIN c1_dbg_r0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END c1_dbg_r0[14]
  PIN c1_dbg_r0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END c1_dbg_r0[15]
  PIN c1_dbg_r0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END c1_dbg_r0[1]
  PIN c1_dbg_r0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END c1_dbg_r0[2]
  PIN c1_dbg_r0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END c1_dbg_r0[3]
  PIN c1_dbg_r0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END c1_dbg_r0[4]
  PIN c1_dbg_r0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END c1_dbg_r0[5]
  PIN c1_dbg_r0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END c1_dbg_r0[6]
  PIN c1_dbg_r0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END c1_dbg_r0[7]
  PIN c1_dbg_r0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END c1_dbg_r0[8]
  PIN c1_dbg_r0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END c1_dbg_r0[9]
  PIN c1_disable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END c1_disable
  PIN c1_i_core_int_sreg[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END c1_i_core_int_sreg[0]
  PIN c1_i_core_int_sreg[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END c1_i_core_int_sreg[10]
  PIN c1_i_core_int_sreg[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END c1_i_core_int_sreg[11]
  PIN c1_i_core_int_sreg[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END c1_i_core_int_sreg[12]
  PIN c1_i_core_int_sreg[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END c1_i_core_int_sreg[13]
  PIN c1_i_core_int_sreg[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END c1_i_core_int_sreg[14]
  PIN c1_i_core_int_sreg[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END c1_i_core_int_sreg[15]
  PIN c1_i_core_int_sreg[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END c1_i_core_int_sreg[1]
  PIN c1_i_core_int_sreg[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END c1_i_core_int_sreg[2]
  PIN c1_i_core_int_sreg[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END c1_i_core_int_sreg[3]
  PIN c1_i_core_int_sreg[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END c1_i_core_int_sreg[4]
  PIN c1_i_core_int_sreg[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END c1_i_core_int_sreg[5]
  PIN c1_i_core_int_sreg[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END c1_i_core_int_sreg[6]
  PIN c1_i_core_int_sreg[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END c1_i_core_int_sreg[7]
  PIN c1_i_core_int_sreg[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 560.360 4.000 560.960 ;
    END
  END c1_i_core_int_sreg[8]
  PIN c1_i_core_int_sreg[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END c1_i_core_int_sreg[9]
  PIN c1_i_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END c1_i_irq
  PIN c1_i_mc_core_int
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END c1_i_mc_core_int
  PIN c1_i_mem_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END c1_i_mem_ack
  PIN c1_i_mem_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END c1_i_mem_data[0]
  PIN c1_i_mem_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END c1_i_mem_data[10]
  PIN c1_i_mem_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END c1_i_mem_data[11]
  PIN c1_i_mem_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END c1_i_mem_data[12]
  PIN c1_i_mem_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END c1_i_mem_data[13]
  PIN c1_i_mem_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END c1_i_mem_data[14]
  PIN c1_i_mem_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.920 4.000 657.520 ;
    END
  END c1_i_mem_data[15]
  PIN c1_i_mem_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END c1_i_mem_data[1]
  PIN c1_i_mem_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END c1_i_mem_data[2]
  PIN c1_i_mem_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END c1_i_mem_data[3]
  PIN c1_i_mem_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END c1_i_mem_data[4]
  PIN c1_i_mem_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END c1_i_mem_data[5]
  PIN c1_i_mem_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END c1_i_mem_data[6]
  PIN c1_i_mem_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END c1_i_mem_data[7]
  PIN c1_i_mem_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END c1_i_mem_data[8]
  PIN c1_i_mem_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END c1_i_mem_data[9]
  PIN c1_i_mem_exception
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END c1_i_mem_exception
  PIN c1_i_req_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END c1_i_req_data[0]
  PIN c1_i_req_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END c1_i_req_data[10]
  PIN c1_i_req_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.880 4.000 604.480 ;
    END
  END c1_i_req_data[11]
  PIN c1_i_req_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END c1_i_req_data[12]
  PIN c1_i_req_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END c1_i_req_data[13]
  PIN c1_i_req_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END c1_i_req_data[14]
  PIN c1_i_req_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END c1_i_req_data[15]
  PIN c1_i_req_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END c1_i_req_data[16]
  PIN c1_i_req_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END c1_i_req_data[17]
  PIN c1_i_req_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END c1_i_req_data[18]
  PIN c1_i_req_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END c1_i_req_data[19]
  PIN c1_i_req_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END c1_i_req_data[1]
  PIN c1_i_req_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END c1_i_req_data[20]
  PIN c1_i_req_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END c1_i_req_data[21]
  PIN c1_i_req_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END c1_i_req_data[22]
  PIN c1_i_req_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END c1_i_req_data[23]
  PIN c1_i_req_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END c1_i_req_data[24]
  PIN c1_i_req_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END c1_i_req_data[25]
  PIN c1_i_req_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END c1_i_req_data[26]
  PIN c1_i_req_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END c1_i_req_data[27]
  PIN c1_i_req_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END c1_i_req_data[28]
  PIN c1_i_req_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END c1_i_req_data[29]
  PIN c1_i_req_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END c1_i_req_data[2]
  PIN c1_i_req_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END c1_i_req_data[30]
  PIN c1_i_req_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END c1_i_req_data[31]
  PIN c1_i_req_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END c1_i_req_data[3]
  PIN c1_i_req_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END c1_i_req_data[4]
  PIN c1_i_req_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END c1_i_req_data[5]
  PIN c1_i_req_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END c1_i_req_data[6]
  PIN c1_i_req_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END c1_i_req_data[7]
  PIN c1_i_req_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END c1_i_req_data[8]
  PIN c1_i_req_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END c1_i_req_data[9]
  PIN c1_i_req_data_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END c1_i_req_data_valid
  PIN c1_o_c_data_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END c1_o_c_data_page
  PIN c1_o_c_instr_long
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END c1_o_c_instr_long
  PIN c1_o_c_instr_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END c1_o_c_instr_page
  PIN c1_o_icache_flush
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END c1_o_icache_flush
  PIN c1_o_instr_long_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END c1_o_instr_long_addr[0]
  PIN c1_o_instr_long_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END c1_o_instr_long_addr[1]
  PIN c1_o_instr_long_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END c1_o_instr_long_addr[2]
  PIN c1_o_instr_long_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END c1_o_instr_long_addr[3]
  PIN c1_o_instr_long_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END c1_o_instr_long_addr[4]
  PIN c1_o_instr_long_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END c1_o_instr_long_addr[5]
  PIN c1_o_instr_long_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END c1_o_instr_long_addr[6]
  PIN c1_o_instr_long_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END c1_o_instr_long_addr[7]
  PIN c1_o_mem_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END c1_o_mem_addr[0]
  PIN c1_o_mem_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END c1_o_mem_addr[10]
  PIN c1_o_mem_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END c1_o_mem_addr[11]
  PIN c1_o_mem_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END c1_o_mem_addr[12]
  PIN c1_o_mem_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END c1_o_mem_addr[13]
  PIN c1_o_mem_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END c1_o_mem_addr[14]
  PIN c1_o_mem_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END c1_o_mem_addr[15]
  PIN c1_o_mem_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END c1_o_mem_addr[1]
  PIN c1_o_mem_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END c1_o_mem_addr[2]
  PIN c1_o_mem_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END c1_o_mem_addr[3]
  PIN c1_o_mem_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END c1_o_mem_addr[4]
  PIN c1_o_mem_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END c1_o_mem_addr[5]
  PIN c1_o_mem_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END c1_o_mem_addr[6]
  PIN c1_o_mem_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END c1_o_mem_addr[7]
  PIN c1_o_mem_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END c1_o_mem_addr[8]
  PIN c1_o_mem_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END c1_o_mem_addr[9]
  PIN c1_o_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END c1_o_mem_data[0]
  PIN c1_o_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END c1_o_mem_data[10]
  PIN c1_o_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END c1_o_mem_data[11]
  PIN c1_o_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END c1_o_mem_data[12]
  PIN c1_o_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END c1_o_mem_data[13]
  PIN c1_o_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END c1_o_mem_data[14]
  PIN c1_o_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END c1_o_mem_data[15]
  PIN c1_o_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END c1_o_mem_data[1]
  PIN c1_o_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END c1_o_mem_data[2]
  PIN c1_o_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END c1_o_mem_data[3]
  PIN c1_o_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END c1_o_mem_data[4]
  PIN c1_o_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END c1_o_mem_data[5]
  PIN c1_o_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END c1_o_mem_data[6]
  PIN c1_o_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END c1_o_mem_data[7]
  PIN c1_o_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END c1_o_mem_data[8]
  PIN c1_o_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END c1_o_mem_data[9]
  PIN c1_o_mem_high_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END c1_o_mem_high_addr[0]
  PIN c1_o_mem_high_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END c1_o_mem_high_addr[1]
  PIN c1_o_mem_high_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END c1_o_mem_high_addr[2]
  PIN c1_o_mem_high_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END c1_o_mem_high_addr[3]
  PIN c1_o_mem_high_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END c1_o_mem_high_addr[4]
  PIN c1_o_mem_high_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END c1_o_mem_high_addr[5]
  PIN c1_o_mem_high_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END c1_o_mem_high_addr[6]
  PIN c1_o_mem_high_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END c1_o_mem_high_addr[7]
  PIN c1_o_mem_long_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END c1_o_mem_long_mode
  PIN c1_o_mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END c1_o_mem_req
  PIN c1_o_mem_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END c1_o_mem_sel[0]
  PIN c1_o_mem_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END c1_o_mem_sel[1]
  PIN c1_o_mem_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END c1_o_mem_we
  PIN c1_o_req_active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END c1_o_req_active
  PIN c1_o_req_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END c1_o_req_addr[0]
  PIN c1_o_req_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END c1_o_req_addr[10]
  PIN c1_o_req_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END c1_o_req_addr[11]
  PIN c1_o_req_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END c1_o_req_addr[12]
  PIN c1_o_req_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END c1_o_req_addr[13]
  PIN c1_o_req_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END c1_o_req_addr[14]
  PIN c1_o_req_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END c1_o_req_addr[15]
  PIN c1_o_req_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END c1_o_req_addr[1]
  PIN c1_o_req_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END c1_o_req_addr[2]
  PIN c1_o_req_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END c1_o_req_addr[3]
  PIN c1_o_req_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END c1_o_req_addr[4]
  PIN c1_o_req_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END c1_o_req_addr[5]
  PIN c1_o_req_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END c1_o_req_addr[6]
  PIN c1_o_req_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END c1_o_req_addr[7]
  PIN c1_o_req_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END c1_o_req_addr[8]
  PIN c1_o_req_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END c1_o_req_addr[9]
  PIN c1_o_req_ppl_submit
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END c1_o_req_ppl_submit
  PIN c1_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END c1_rst
  PIN c1_sr_bus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END c1_sr_bus_addr[0]
  PIN c1_sr_bus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END c1_sr_bus_addr[10]
  PIN c1_sr_bus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END c1_sr_bus_addr[11]
  PIN c1_sr_bus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END c1_sr_bus_addr[12]
  PIN c1_sr_bus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END c1_sr_bus_addr[13]
  PIN c1_sr_bus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END c1_sr_bus_addr[14]
  PIN c1_sr_bus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.720 4.000 664.320 ;
    END
  END c1_sr_bus_addr[15]
  PIN c1_sr_bus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END c1_sr_bus_addr[1]
  PIN c1_sr_bus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END c1_sr_bus_addr[2]
  PIN c1_sr_bus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END c1_sr_bus_addr[3]
  PIN c1_sr_bus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END c1_sr_bus_addr[4]
  PIN c1_sr_bus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END c1_sr_bus_addr[5]
  PIN c1_sr_bus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END c1_sr_bus_addr[6]
  PIN c1_sr_bus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END c1_sr_bus_addr[7]
  PIN c1_sr_bus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END c1_sr_bus_addr[8]
  PIN c1_sr_bus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END c1_sr_bus_addr[9]
  PIN c1_sr_bus_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END c1_sr_bus_data_o[0]
  PIN c1_sr_bus_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END c1_sr_bus_data_o[10]
  PIN c1_sr_bus_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END c1_sr_bus_data_o[11]
  PIN c1_sr_bus_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END c1_sr_bus_data_o[12]
  PIN c1_sr_bus_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END c1_sr_bus_data_o[13]
  PIN c1_sr_bus_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 651.480 4.000 652.080 ;
    END
  END c1_sr_bus_data_o[14]
  PIN c1_sr_bus_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END c1_sr_bus_data_o[15]
  PIN c1_sr_bus_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END c1_sr_bus_data_o[1]
  PIN c1_sr_bus_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END c1_sr_bus_data_o[2]
  PIN c1_sr_bus_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END c1_sr_bus_data_o[3]
  PIN c1_sr_bus_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END c1_sr_bus_data_o[4]
  PIN c1_sr_bus_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END c1_sr_bus_data_o[5]
  PIN c1_sr_bus_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END c1_sr_bus_data_o[6]
  PIN c1_sr_bus_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END c1_sr_bus_data_o[7]
  PIN c1_sr_bus_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END c1_sr_bus_data_o[8]
  PIN c1_sr_bus_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END c1_sr_bus_data_o[9]
  PIN c1_sr_bus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END c1_sr_bus_we
  PIN core_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END core_clock
  PIN core_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END core_reset
  PIN dcache_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 78.920 300.000 79.520 ;
    END
  END dcache_clk
  PIN dcache_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 80.960 300.000 81.560 ;
    END
  END dcache_mem_ack
  PIN dcache_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 105.440 300.000 106.040 ;
    END
  END dcache_mem_addr[0]
  PIN dcache_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 236.000 300.000 236.600 ;
    END
  END dcache_mem_addr[10]
  PIN dcache_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 248.240 300.000 248.840 ;
    END
  END dcache_mem_addr[11]
  PIN dcache_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 260.480 300.000 261.080 ;
    END
  END dcache_mem_addr[12]
  PIN dcache_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 272.720 300.000 273.320 ;
    END
  END dcache_mem_addr[13]
  PIN dcache_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 284.960 300.000 285.560 ;
    END
  END dcache_mem_addr[14]
  PIN dcache_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 297.200 300.000 297.800 ;
    END
  END dcache_mem_addr[15]
  PIN dcache_mem_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 309.440 300.000 310.040 ;
    END
  END dcache_mem_addr[16]
  PIN dcache_mem_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 313.520 300.000 314.120 ;
    END
  END dcache_mem_addr[17]
  PIN dcache_mem_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 317.600 300.000 318.200 ;
    END
  END dcache_mem_addr[18]
  PIN dcache_mem_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 321.680 300.000 322.280 ;
    END
  END dcache_mem_addr[19]
  PIN dcache_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 121.760 300.000 122.360 ;
    END
  END dcache_mem_addr[1]
  PIN dcache_mem_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 325.760 300.000 326.360 ;
    END
  END dcache_mem_addr[20]
  PIN dcache_mem_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 329.840 300.000 330.440 ;
    END
  END dcache_mem_addr[21]
  PIN dcache_mem_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 333.920 300.000 334.520 ;
    END
  END dcache_mem_addr[22]
  PIN dcache_mem_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 338.000 300.000 338.600 ;
    END
  END dcache_mem_addr[23]
  PIN dcache_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 138.080 300.000 138.680 ;
    END
  END dcache_mem_addr[2]
  PIN dcache_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 150.320 300.000 150.920 ;
    END
  END dcache_mem_addr[3]
  PIN dcache_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 162.560 300.000 163.160 ;
    END
  END dcache_mem_addr[4]
  PIN dcache_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 174.800 300.000 175.400 ;
    END
  END dcache_mem_addr[5]
  PIN dcache_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 187.040 300.000 187.640 ;
    END
  END dcache_mem_addr[6]
  PIN dcache_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 199.280 300.000 199.880 ;
    END
  END dcache_mem_addr[7]
  PIN dcache_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 211.520 300.000 212.120 ;
    END
  END dcache_mem_addr[8]
  PIN dcache_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 223.760 300.000 224.360 ;
    END
  END dcache_mem_addr[9]
  PIN dcache_mem_cache_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 83.000 300.000 83.600 ;
    END
  END dcache_mem_cache_enable
  PIN dcache_mem_exception
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 85.040 300.000 85.640 ;
    END
  END dcache_mem_exception
  PIN dcache_mem_i_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.480 300.000 108.080 ;
    END
  END dcache_mem_i_data[0]
  PIN dcache_mem_i_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 238.040 300.000 238.640 ;
    END
  END dcache_mem_i_data[10]
  PIN dcache_mem_i_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 250.280 300.000 250.880 ;
    END
  END dcache_mem_i_data[11]
  PIN dcache_mem_i_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 262.520 300.000 263.120 ;
    END
  END dcache_mem_i_data[12]
  PIN dcache_mem_i_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 274.760 300.000 275.360 ;
    END
  END dcache_mem_i_data[13]
  PIN dcache_mem_i_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 287.000 300.000 287.600 ;
    END
  END dcache_mem_i_data[14]
  PIN dcache_mem_i_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 299.240 300.000 299.840 ;
    END
  END dcache_mem_i_data[15]
  PIN dcache_mem_i_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 123.800 300.000 124.400 ;
    END
  END dcache_mem_i_data[1]
  PIN dcache_mem_i_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 140.120 300.000 140.720 ;
    END
  END dcache_mem_i_data[2]
  PIN dcache_mem_i_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 152.360 300.000 152.960 ;
    END
  END dcache_mem_i_data[3]
  PIN dcache_mem_i_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.600 300.000 165.200 ;
    END
  END dcache_mem_i_data[4]
  PIN dcache_mem_i_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.840 300.000 177.440 ;
    END
  END dcache_mem_i_data[5]
  PIN dcache_mem_i_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 189.080 300.000 189.680 ;
    END
  END dcache_mem_i_data[6]
  PIN dcache_mem_i_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.320 300.000 201.920 ;
    END
  END dcache_mem_i_data[7]
  PIN dcache_mem_i_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 213.560 300.000 214.160 ;
    END
  END dcache_mem_i_data[8]
  PIN dcache_mem_i_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 225.800 300.000 226.400 ;
    END
  END dcache_mem_i_data[9]
  PIN dcache_mem_o_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 109.520 300.000 110.120 ;
    END
  END dcache_mem_o_data[0]
  PIN dcache_mem_o_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 240.080 300.000 240.680 ;
    END
  END dcache_mem_o_data[10]
  PIN dcache_mem_o_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 252.320 300.000 252.920 ;
    END
  END dcache_mem_o_data[11]
  PIN dcache_mem_o_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 264.560 300.000 265.160 ;
    END
  END dcache_mem_o_data[12]
  PIN dcache_mem_o_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 276.800 300.000 277.400 ;
    END
  END dcache_mem_o_data[13]
  PIN dcache_mem_o_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.040 300.000 289.640 ;
    END
  END dcache_mem_o_data[14]
  PIN dcache_mem_o_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 301.280 300.000 301.880 ;
    END
  END dcache_mem_o_data[15]
  PIN dcache_mem_o_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.840 300.000 126.440 ;
    END
  END dcache_mem_o_data[1]
  PIN dcache_mem_o_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 142.160 300.000 142.760 ;
    END
  END dcache_mem_o_data[2]
  PIN dcache_mem_o_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 154.400 300.000 155.000 ;
    END
  END dcache_mem_o_data[3]
  PIN dcache_mem_o_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 166.640 300.000 167.240 ;
    END
  END dcache_mem_o_data[4]
  PIN dcache_mem_o_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 178.880 300.000 179.480 ;
    END
  END dcache_mem_o_data[5]
  PIN dcache_mem_o_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 191.120 300.000 191.720 ;
    END
  END dcache_mem_o_data[6]
  PIN dcache_mem_o_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 203.360 300.000 203.960 ;
    END
  END dcache_mem_o_data[7]
  PIN dcache_mem_o_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 215.600 300.000 216.200 ;
    END
  END dcache_mem_o_data[8]
  PIN dcache_mem_o_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 227.840 300.000 228.440 ;
    END
  END dcache_mem_o_data[9]
  PIN dcache_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 87.080 300.000 87.680 ;
    END
  END dcache_mem_req
  PIN dcache_mem_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.560 300.000 112.160 ;
    END
  END dcache_mem_sel[0]
  PIN dcache_mem_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 127.880 300.000 128.480 ;
    END
  END dcache_mem_sel[1]
  PIN dcache_mem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 89.120 300.000 89.720 ;
    END
  END dcache_mem_we
  PIN dcache_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.160 300.000 91.760 ;
    END
  END dcache_rst
  PIN dcache_wb_4_burst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 93.200 300.000 93.800 ;
    END
  END dcache_wb_4_burst
  PIN dcache_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 95.240 300.000 95.840 ;
    END
  END dcache_wb_ack
  PIN dcache_wb_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 113.600 300.000 114.200 ;
    END
  END dcache_wb_adr[0]
  PIN dcache_wb_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 242.120 300.000 242.720 ;
    END
  END dcache_wb_adr[10]
  PIN dcache_wb_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 254.360 300.000 254.960 ;
    END
  END dcache_wb_adr[11]
  PIN dcache_wb_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.600 300.000 267.200 ;
    END
  END dcache_wb_adr[12]
  PIN dcache_wb_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 278.840 300.000 279.440 ;
    END
  END dcache_wb_adr[13]
  PIN dcache_wb_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 291.080 300.000 291.680 ;
    END
  END dcache_wb_adr[14]
  PIN dcache_wb_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 303.320 300.000 303.920 ;
    END
  END dcache_wb_adr[15]
  PIN dcache_wb_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 311.480 300.000 312.080 ;
    END
  END dcache_wb_adr[16]
  PIN dcache_wb_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 315.560 300.000 316.160 ;
    END
  END dcache_wb_adr[17]
  PIN dcache_wb_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 319.640 300.000 320.240 ;
    END
  END dcache_wb_adr[18]
  PIN dcache_wb_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 323.720 300.000 324.320 ;
    END
  END dcache_wb_adr[19]
  PIN dcache_wb_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 129.920 300.000 130.520 ;
    END
  END dcache_wb_adr[1]
  PIN dcache_wb_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 327.800 300.000 328.400 ;
    END
  END dcache_wb_adr[20]
  PIN dcache_wb_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 331.880 300.000 332.480 ;
    END
  END dcache_wb_adr[21]
  PIN dcache_wb_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 335.960 300.000 336.560 ;
    END
  END dcache_wb_adr[22]
  PIN dcache_wb_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 340.040 300.000 340.640 ;
    END
  END dcache_wb_adr[23]
  PIN dcache_wb_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 144.200 300.000 144.800 ;
    END
  END dcache_wb_adr[2]
  PIN dcache_wb_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.440 300.000 157.040 ;
    END
  END dcache_wb_adr[3]
  PIN dcache_wb_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 168.680 300.000 169.280 ;
    END
  END dcache_wb_adr[4]
  PIN dcache_wb_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 180.920 300.000 181.520 ;
    END
  END dcache_wb_adr[5]
  PIN dcache_wb_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 193.160 300.000 193.760 ;
    END
  END dcache_wb_adr[6]
  PIN dcache_wb_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.400 300.000 206.000 ;
    END
  END dcache_wb_adr[7]
  PIN dcache_wb_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 217.640 300.000 218.240 ;
    END
  END dcache_wb_adr[8]
  PIN dcache_wb_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 229.880 300.000 230.480 ;
    END
  END dcache_wb_adr[9]
  PIN dcache_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 97.280 300.000 97.880 ;
    END
  END dcache_wb_cyc
  PIN dcache_wb_err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 99.320 300.000 99.920 ;
    END
  END dcache_wb_err
  PIN dcache_wb_i_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 115.640 300.000 116.240 ;
    END
  END dcache_wb_i_dat[0]
  PIN dcache_wb_i_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.160 300.000 244.760 ;
    END
  END dcache_wb_i_dat[10]
  PIN dcache_wb_i_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 256.400 300.000 257.000 ;
    END
  END dcache_wb_i_dat[11]
  PIN dcache_wb_i_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.640 300.000 269.240 ;
    END
  END dcache_wb_i_dat[12]
  PIN dcache_wb_i_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 280.880 300.000 281.480 ;
    END
  END dcache_wb_i_dat[13]
  PIN dcache_wb_i_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 293.120 300.000 293.720 ;
    END
  END dcache_wb_i_dat[14]
  PIN dcache_wb_i_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 305.360 300.000 305.960 ;
    END
  END dcache_wb_i_dat[15]
  PIN dcache_wb_i_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 131.960 300.000 132.560 ;
    END
  END dcache_wb_i_dat[1]
  PIN dcache_wb_i_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.240 300.000 146.840 ;
    END
  END dcache_wb_i_dat[2]
  PIN dcache_wb_i_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 158.480 300.000 159.080 ;
    END
  END dcache_wb_i_dat[3]
  PIN dcache_wb_i_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 170.720 300.000 171.320 ;
    END
  END dcache_wb_i_dat[4]
  PIN dcache_wb_i_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.960 300.000 183.560 ;
    END
  END dcache_wb_i_dat[5]
  PIN dcache_wb_i_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 195.200 300.000 195.800 ;
    END
  END dcache_wb_i_dat[6]
  PIN dcache_wb_i_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 207.440 300.000 208.040 ;
    END
  END dcache_wb_i_dat[7]
  PIN dcache_wb_i_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 219.680 300.000 220.280 ;
    END
  END dcache_wb_i_dat[8]
  PIN dcache_wb_i_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 231.920 300.000 232.520 ;
    END
  END dcache_wb_i_dat[9]
  PIN dcache_wb_o_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 117.680 300.000 118.280 ;
    END
  END dcache_wb_o_dat[0]
  PIN dcache_wb_o_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 246.200 300.000 246.800 ;
    END
  END dcache_wb_o_dat[10]
  PIN dcache_wb_o_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.440 300.000 259.040 ;
    END
  END dcache_wb_o_dat[11]
  PIN dcache_wb_o_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 270.680 300.000 271.280 ;
    END
  END dcache_wb_o_dat[12]
  PIN dcache_wb_o_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 282.920 300.000 283.520 ;
    END
  END dcache_wb_o_dat[13]
  PIN dcache_wb_o_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 295.160 300.000 295.760 ;
    END
  END dcache_wb_o_dat[14]
  PIN dcache_wb_o_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 307.400 300.000 308.000 ;
    END
  END dcache_wb_o_dat[15]
  PIN dcache_wb_o_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 134.000 300.000 134.600 ;
    END
  END dcache_wb_o_dat[1]
  PIN dcache_wb_o_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.280 300.000 148.880 ;
    END
  END dcache_wb_o_dat[2]
  PIN dcache_wb_o_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 160.520 300.000 161.120 ;
    END
  END dcache_wb_o_dat[3]
  PIN dcache_wb_o_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 172.760 300.000 173.360 ;
    END
  END dcache_wb_o_dat[4]
  PIN dcache_wb_o_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 185.000 300.000 185.600 ;
    END
  END dcache_wb_o_dat[5]
  PIN dcache_wb_o_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 197.240 300.000 197.840 ;
    END
  END dcache_wb_o_dat[6]
  PIN dcache_wb_o_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 209.480 300.000 210.080 ;
    END
  END dcache_wb_o_dat[7]
  PIN dcache_wb_o_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.720 300.000 222.320 ;
    END
  END dcache_wb_o_dat[8]
  PIN dcache_wb_o_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 233.960 300.000 234.560 ;
    END
  END dcache_wb_o_dat[9]
  PIN dcache_wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 119.720 300.000 120.320 ;
    END
  END dcache_wb_sel[0]
  PIN dcache_wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.040 300.000 136.640 ;
    END
  END dcache_wb_sel[1]
  PIN dcache_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 101.360 300.000 101.960 ;
    END
  END dcache_wb_stb
  PIN dcache_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 103.400 300.000 104.000 ;
    END
  END dcache_wb_we
  PIN ic0_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 342.080 300.000 342.680 ;
    END
  END ic0_clk
  PIN ic0_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 344.120 300.000 344.720 ;
    END
  END ic0_mem_ack
  PIN ic0_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 364.520 300.000 365.120 ;
    END
  END ic0_mem_addr[0]
  PIN ic0_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 450.200 300.000 450.800 ;
    END
  END ic0_mem_addr[10]
  PIN ic0_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 458.360 300.000 458.960 ;
    END
  END ic0_mem_addr[11]
  PIN ic0_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 466.520 300.000 467.120 ;
    END
  END ic0_mem_addr[12]
  PIN ic0_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 474.680 300.000 475.280 ;
    END
  END ic0_mem_addr[13]
  PIN ic0_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 482.840 300.000 483.440 ;
    END
  END ic0_mem_addr[14]
  PIN ic0_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 491.000 300.000 491.600 ;
    END
  END ic0_mem_addr[15]
  PIN ic0_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 374.720 300.000 375.320 ;
    END
  END ic0_mem_addr[1]
  PIN ic0_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 384.920 300.000 385.520 ;
    END
  END ic0_mem_addr[2]
  PIN ic0_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 393.080 300.000 393.680 ;
    END
  END ic0_mem_addr[3]
  PIN ic0_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 401.240 300.000 401.840 ;
    END
  END ic0_mem_addr[4]
  PIN ic0_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 409.400 300.000 410.000 ;
    END
  END ic0_mem_addr[5]
  PIN ic0_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 417.560 300.000 418.160 ;
    END
  END ic0_mem_addr[6]
  PIN ic0_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 425.720 300.000 426.320 ;
    END
  END ic0_mem_addr[7]
  PIN ic0_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 433.880 300.000 434.480 ;
    END
  END ic0_mem_addr[8]
  PIN ic0_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 442.040 300.000 442.640 ;
    END
  END ic0_mem_addr[9]
  PIN ic0_mem_cache_flush
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 346.160 300.000 346.760 ;
    END
  END ic0_mem_cache_flush
  PIN ic0_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 366.560 300.000 367.160 ;
    END
  END ic0_mem_data[0]
  PIN ic0_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 452.240 300.000 452.840 ;
    END
  END ic0_mem_data[10]
  PIN ic0_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 460.400 300.000 461.000 ;
    END
  END ic0_mem_data[11]
  PIN ic0_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 468.560 300.000 469.160 ;
    END
  END ic0_mem_data[12]
  PIN ic0_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 476.720 300.000 477.320 ;
    END
  END ic0_mem_data[13]
  PIN ic0_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 484.880 300.000 485.480 ;
    END
  END ic0_mem_data[14]
  PIN ic0_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 493.040 300.000 493.640 ;
    END
  END ic0_mem_data[15]
  PIN ic0_mem_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 499.160 300.000 499.760 ;
    END
  END ic0_mem_data[16]
  PIN ic0_mem_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 501.200 300.000 501.800 ;
    END
  END ic0_mem_data[17]
  PIN ic0_mem_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 503.240 300.000 503.840 ;
    END
  END ic0_mem_data[18]
  PIN ic0_mem_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 505.280 300.000 505.880 ;
    END
  END ic0_mem_data[19]
  PIN ic0_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 376.760 300.000 377.360 ;
    END
  END ic0_mem_data[1]
  PIN ic0_mem_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 507.320 300.000 507.920 ;
    END
  END ic0_mem_data[20]
  PIN ic0_mem_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 509.360 300.000 509.960 ;
    END
  END ic0_mem_data[21]
  PIN ic0_mem_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 511.400 300.000 512.000 ;
    END
  END ic0_mem_data[22]
  PIN ic0_mem_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 513.440 300.000 514.040 ;
    END
  END ic0_mem_data[23]
  PIN ic0_mem_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 515.480 300.000 516.080 ;
    END
  END ic0_mem_data[24]
  PIN ic0_mem_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 517.520 300.000 518.120 ;
    END
  END ic0_mem_data[25]
  PIN ic0_mem_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 519.560 300.000 520.160 ;
    END
  END ic0_mem_data[26]
  PIN ic0_mem_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 521.600 300.000 522.200 ;
    END
  END ic0_mem_data[27]
  PIN ic0_mem_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 523.640 300.000 524.240 ;
    END
  END ic0_mem_data[28]
  PIN ic0_mem_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 525.680 300.000 526.280 ;
    END
  END ic0_mem_data[29]
  PIN ic0_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 386.960 300.000 387.560 ;
    END
  END ic0_mem_data[2]
  PIN ic0_mem_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 527.720 300.000 528.320 ;
    END
  END ic0_mem_data[30]
  PIN ic0_mem_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 529.760 300.000 530.360 ;
    END
  END ic0_mem_data[31]
  PIN ic0_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 395.120 300.000 395.720 ;
    END
  END ic0_mem_data[3]
  PIN ic0_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 403.280 300.000 403.880 ;
    END
  END ic0_mem_data[4]
  PIN ic0_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 411.440 300.000 412.040 ;
    END
  END ic0_mem_data[5]
  PIN ic0_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 419.600 300.000 420.200 ;
    END
  END ic0_mem_data[6]
  PIN ic0_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 427.760 300.000 428.360 ;
    END
  END ic0_mem_data[7]
  PIN ic0_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 435.920 300.000 436.520 ;
    END
  END ic0_mem_data[8]
  PIN ic0_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 444.080 300.000 444.680 ;
    END
  END ic0_mem_data[9]
  PIN ic0_mem_ppl_submit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 348.200 300.000 348.800 ;
    END
  END ic0_mem_ppl_submit
  PIN ic0_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 350.240 300.000 350.840 ;
    END
  END ic0_mem_req
  PIN ic0_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 352.280 300.000 352.880 ;
    END
  END ic0_rst
  PIN ic0_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 354.320 300.000 354.920 ;
    END
  END ic0_wb_ack
  PIN ic0_wb_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 368.600 300.000 369.200 ;
    END
  END ic0_wb_adr[0]
  PIN ic0_wb_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 454.280 300.000 454.880 ;
    END
  END ic0_wb_adr[10]
  PIN ic0_wb_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 462.440 300.000 463.040 ;
    END
  END ic0_wb_adr[11]
  PIN ic0_wb_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 470.600 300.000 471.200 ;
    END
  END ic0_wb_adr[12]
  PIN ic0_wb_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 478.760 300.000 479.360 ;
    END
  END ic0_wb_adr[13]
  PIN ic0_wb_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 486.920 300.000 487.520 ;
    END
  END ic0_wb_adr[14]
  PIN ic0_wb_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 495.080 300.000 495.680 ;
    END
  END ic0_wb_adr[15]
  PIN ic0_wb_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 378.800 300.000 379.400 ;
    END
  END ic0_wb_adr[1]
  PIN ic0_wb_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 389.000 300.000 389.600 ;
    END
  END ic0_wb_adr[2]
  PIN ic0_wb_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 397.160 300.000 397.760 ;
    END
  END ic0_wb_adr[3]
  PIN ic0_wb_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 405.320 300.000 405.920 ;
    END
  END ic0_wb_adr[4]
  PIN ic0_wb_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 413.480 300.000 414.080 ;
    END
  END ic0_wb_adr[5]
  PIN ic0_wb_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 421.640 300.000 422.240 ;
    END
  END ic0_wb_adr[6]
  PIN ic0_wb_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 429.800 300.000 430.400 ;
    END
  END ic0_wb_adr[7]
  PIN ic0_wb_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 437.960 300.000 438.560 ;
    END
  END ic0_wb_adr[8]
  PIN ic0_wb_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 446.120 300.000 446.720 ;
    END
  END ic0_wb_adr[9]
  PIN ic0_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 356.360 300.000 356.960 ;
    END
  END ic0_wb_cyc
  PIN ic0_wb_err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 358.400 300.000 359.000 ;
    END
  END ic0_wb_err
  PIN ic0_wb_i_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 370.640 300.000 371.240 ;
    END
  END ic0_wb_i_dat[0]
  PIN ic0_wb_i_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 456.320 300.000 456.920 ;
    END
  END ic0_wb_i_dat[10]
  PIN ic0_wb_i_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 464.480 300.000 465.080 ;
    END
  END ic0_wb_i_dat[11]
  PIN ic0_wb_i_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 472.640 300.000 473.240 ;
    END
  END ic0_wb_i_dat[12]
  PIN ic0_wb_i_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 480.800 300.000 481.400 ;
    END
  END ic0_wb_i_dat[13]
  PIN ic0_wb_i_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 488.960 300.000 489.560 ;
    END
  END ic0_wb_i_dat[14]
  PIN ic0_wb_i_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 497.120 300.000 497.720 ;
    END
  END ic0_wb_i_dat[15]
  PIN ic0_wb_i_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 380.840 300.000 381.440 ;
    END
  END ic0_wb_i_dat[1]
  PIN ic0_wb_i_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 391.040 300.000 391.640 ;
    END
  END ic0_wb_i_dat[2]
  PIN ic0_wb_i_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 399.200 300.000 399.800 ;
    END
  END ic0_wb_i_dat[3]
  PIN ic0_wb_i_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 407.360 300.000 407.960 ;
    END
  END ic0_wb_i_dat[4]
  PIN ic0_wb_i_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 415.520 300.000 416.120 ;
    END
  END ic0_wb_i_dat[5]
  PIN ic0_wb_i_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 423.680 300.000 424.280 ;
    END
  END ic0_wb_i_dat[6]
  PIN ic0_wb_i_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 431.840 300.000 432.440 ;
    END
  END ic0_wb_i_dat[7]
  PIN ic0_wb_i_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 440.000 300.000 440.600 ;
    END
  END ic0_wb_i_dat[8]
  PIN ic0_wb_i_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 448.160 300.000 448.760 ;
    END
  END ic0_wb_i_dat[9]
  PIN ic0_wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 372.680 300.000 373.280 ;
    END
  END ic0_wb_sel[0]
  PIN ic0_wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 382.880 300.000 383.480 ;
    END
  END ic0_wb_sel[1]
  PIN ic0_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 360.440 300.000 361.040 ;
    END
  END ic0_wb_stb
  PIN ic0_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 362.480 300.000 363.080 ;
    END
  END ic0_wb_we
  PIN ic1_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 531.800 300.000 532.400 ;
    END
  END ic1_clk
  PIN ic1_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 533.840 300.000 534.440 ;
    END
  END ic1_mem_ack
  PIN ic1_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 554.240 300.000 554.840 ;
    END
  END ic1_mem_addr[0]
  PIN ic1_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 639.920 300.000 640.520 ;
    END
  END ic1_mem_addr[10]
  PIN ic1_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 648.080 300.000 648.680 ;
    END
  END ic1_mem_addr[11]
  PIN ic1_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 656.240 300.000 656.840 ;
    END
  END ic1_mem_addr[12]
  PIN ic1_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 664.400 300.000 665.000 ;
    END
  END ic1_mem_addr[13]
  PIN ic1_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 672.560 300.000 673.160 ;
    END
  END ic1_mem_addr[14]
  PIN ic1_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 680.720 300.000 681.320 ;
    END
  END ic1_mem_addr[15]
  PIN ic1_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 564.440 300.000 565.040 ;
    END
  END ic1_mem_addr[1]
  PIN ic1_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 574.640 300.000 575.240 ;
    END
  END ic1_mem_addr[2]
  PIN ic1_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 582.800 300.000 583.400 ;
    END
  END ic1_mem_addr[3]
  PIN ic1_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 590.960 300.000 591.560 ;
    END
  END ic1_mem_addr[4]
  PIN ic1_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 599.120 300.000 599.720 ;
    END
  END ic1_mem_addr[5]
  PIN ic1_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 607.280 300.000 607.880 ;
    END
  END ic1_mem_addr[6]
  PIN ic1_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 615.440 300.000 616.040 ;
    END
  END ic1_mem_addr[7]
  PIN ic1_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 623.600 300.000 624.200 ;
    END
  END ic1_mem_addr[8]
  PIN ic1_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 631.760 300.000 632.360 ;
    END
  END ic1_mem_addr[9]
  PIN ic1_mem_cache_flush
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 535.880 300.000 536.480 ;
    END
  END ic1_mem_cache_flush
  PIN ic1_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 556.280 300.000 556.880 ;
    END
  END ic1_mem_data[0]
  PIN ic1_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 641.960 300.000 642.560 ;
    END
  END ic1_mem_data[10]
  PIN ic1_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 650.120 300.000 650.720 ;
    END
  END ic1_mem_data[11]
  PIN ic1_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 658.280 300.000 658.880 ;
    END
  END ic1_mem_data[12]
  PIN ic1_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 666.440 300.000 667.040 ;
    END
  END ic1_mem_data[13]
  PIN ic1_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 674.600 300.000 675.200 ;
    END
  END ic1_mem_data[14]
  PIN ic1_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 682.760 300.000 683.360 ;
    END
  END ic1_mem_data[15]
  PIN ic1_mem_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 688.880 300.000 689.480 ;
    END
  END ic1_mem_data[16]
  PIN ic1_mem_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 690.920 300.000 691.520 ;
    END
  END ic1_mem_data[17]
  PIN ic1_mem_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 692.960 300.000 693.560 ;
    END
  END ic1_mem_data[18]
  PIN ic1_mem_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 695.000 300.000 695.600 ;
    END
  END ic1_mem_data[19]
  PIN ic1_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 566.480 300.000 567.080 ;
    END
  END ic1_mem_data[1]
  PIN ic1_mem_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 697.040 300.000 697.640 ;
    END
  END ic1_mem_data[20]
  PIN ic1_mem_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 699.080 300.000 699.680 ;
    END
  END ic1_mem_data[21]
  PIN ic1_mem_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 701.120 300.000 701.720 ;
    END
  END ic1_mem_data[22]
  PIN ic1_mem_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 703.160 300.000 703.760 ;
    END
  END ic1_mem_data[23]
  PIN ic1_mem_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 705.200 300.000 705.800 ;
    END
  END ic1_mem_data[24]
  PIN ic1_mem_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 707.240 300.000 707.840 ;
    END
  END ic1_mem_data[25]
  PIN ic1_mem_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 709.280 300.000 709.880 ;
    END
  END ic1_mem_data[26]
  PIN ic1_mem_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 711.320 300.000 711.920 ;
    END
  END ic1_mem_data[27]
  PIN ic1_mem_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 713.360 300.000 713.960 ;
    END
  END ic1_mem_data[28]
  PIN ic1_mem_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 715.400 300.000 716.000 ;
    END
  END ic1_mem_data[29]
  PIN ic1_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 576.680 300.000 577.280 ;
    END
  END ic1_mem_data[2]
  PIN ic1_mem_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 717.440 300.000 718.040 ;
    END
  END ic1_mem_data[30]
  PIN ic1_mem_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 719.480 300.000 720.080 ;
    END
  END ic1_mem_data[31]
  PIN ic1_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 584.840 300.000 585.440 ;
    END
  END ic1_mem_data[3]
  PIN ic1_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 593.000 300.000 593.600 ;
    END
  END ic1_mem_data[4]
  PIN ic1_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 601.160 300.000 601.760 ;
    END
  END ic1_mem_data[5]
  PIN ic1_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 609.320 300.000 609.920 ;
    END
  END ic1_mem_data[6]
  PIN ic1_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 617.480 300.000 618.080 ;
    END
  END ic1_mem_data[7]
  PIN ic1_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 625.640 300.000 626.240 ;
    END
  END ic1_mem_data[8]
  PIN ic1_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 633.800 300.000 634.400 ;
    END
  END ic1_mem_data[9]
  PIN ic1_mem_ppl_submit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 537.920 300.000 538.520 ;
    END
  END ic1_mem_ppl_submit
  PIN ic1_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 539.960 300.000 540.560 ;
    END
  END ic1_mem_req
  PIN ic1_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 542.000 300.000 542.600 ;
    END
  END ic1_rst
  PIN ic1_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 544.040 300.000 544.640 ;
    END
  END ic1_wb_ack
  PIN ic1_wb_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 558.320 300.000 558.920 ;
    END
  END ic1_wb_adr[0]
  PIN ic1_wb_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 644.000 300.000 644.600 ;
    END
  END ic1_wb_adr[10]
  PIN ic1_wb_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 652.160 300.000 652.760 ;
    END
  END ic1_wb_adr[11]
  PIN ic1_wb_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 660.320 300.000 660.920 ;
    END
  END ic1_wb_adr[12]
  PIN ic1_wb_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 668.480 300.000 669.080 ;
    END
  END ic1_wb_adr[13]
  PIN ic1_wb_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 676.640 300.000 677.240 ;
    END
  END ic1_wb_adr[14]
  PIN ic1_wb_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 684.800 300.000 685.400 ;
    END
  END ic1_wb_adr[15]
  PIN ic1_wb_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 568.520 300.000 569.120 ;
    END
  END ic1_wb_adr[1]
  PIN ic1_wb_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 578.720 300.000 579.320 ;
    END
  END ic1_wb_adr[2]
  PIN ic1_wb_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 586.880 300.000 587.480 ;
    END
  END ic1_wb_adr[3]
  PIN ic1_wb_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 595.040 300.000 595.640 ;
    END
  END ic1_wb_adr[4]
  PIN ic1_wb_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 603.200 300.000 603.800 ;
    END
  END ic1_wb_adr[5]
  PIN ic1_wb_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 611.360 300.000 611.960 ;
    END
  END ic1_wb_adr[6]
  PIN ic1_wb_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 619.520 300.000 620.120 ;
    END
  END ic1_wb_adr[7]
  PIN ic1_wb_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 627.680 300.000 628.280 ;
    END
  END ic1_wb_adr[8]
  PIN ic1_wb_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 635.840 300.000 636.440 ;
    END
  END ic1_wb_adr[9]
  PIN ic1_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 546.080 300.000 546.680 ;
    END
  END ic1_wb_cyc
  PIN ic1_wb_err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 548.120 300.000 548.720 ;
    END
  END ic1_wb_err
  PIN ic1_wb_i_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 560.360 300.000 560.960 ;
    END
  END ic1_wb_i_dat[0]
  PIN ic1_wb_i_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 646.040 300.000 646.640 ;
    END
  END ic1_wb_i_dat[10]
  PIN ic1_wb_i_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 654.200 300.000 654.800 ;
    END
  END ic1_wb_i_dat[11]
  PIN ic1_wb_i_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 662.360 300.000 662.960 ;
    END
  END ic1_wb_i_dat[12]
  PIN ic1_wb_i_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 670.520 300.000 671.120 ;
    END
  END ic1_wb_i_dat[13]
  PIN ic1_wb_i_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 678.680 300.000 679.280 ;
    END
  END ic1_wb_i_dat[14]
  PIN ic1_wb_i_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 686.840 300.000 687.440 ;
    END
  END ic1_wb_i_dat[15]
  PIN ic1_wb_i_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 570.560 300.000 571.160 ;
    END
  END ic1_wb_i_dat[1]
  PIN ic1_wb_i_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 580.760 300.000 581.360 ;
    END
  END ic1_wb_i_dat[2]
  PIN ic1_wb_i_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 588.920 300.000 589.520 ;
    END
  END ic1_wb_i_dat[3]
  PIN ic1_wb_i_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 597.080 300.000 597.680 ;
    END
  END ic1_wb_i_dat[4]
  PIN ic1_wb_i_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 605.240 300.000 605.840 ;
    END
  END ic1_wb_i_dat[5]
  PIN ic1_wb_i_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 613.400 300.000 614.000 ;
    END
  END ic1_wb_i_dat[6]
  PIN ic1_wb_i_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 621.560 300.000 622.160 ;
    END
  END ic1_wb_i_dat[7]
  PIN ic1_wb_i_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 629.720 300.000 630.320 ;
    END
  END ic1_wb_i_dat[8]
  PIN ic1_wb_i_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 637.880 300.000 638.480 ;
    END
  END ic1_wb_i_dat[9]
  PIN ic1_wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 562.400 300.000 563.000 ;
    END
  END ic1_wb_sel[0]
  PIN ic1_wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 572.600 300.000 573.200 ;
    END
  END ic1_wb_sel[1]
  PIN ic1_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 550.160 300.000 550.760 ;
    END
  END ic1_wb_stb
  PIN ic1_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 552.200 300.000 552.800 ;
    END
  END ic1_wb_we
  PIN inner_disable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END inner_disable
  PIN inner_embed_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END inner_embed_mode
  PIN inner_ext_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END inner_ext_irq
  PIN inner_wb_4_burst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END inner_wb_4_burst
  PIN inner_wb_8_burst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END inner_wb_8_burst
  PIN inner_wb_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END inner_wb_ack
  PIN inner_wb_adr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END inner_wb_adr[0]
  PIN inner_wb_adr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END inner_wb_adr[10]
  PIN inner_wb_adr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END inner_wb_adr[11]
  PIN inner_wb_adr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END inner_wb_adr[12]
  PIN inner_wb_adr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END inner_wb_adr[13]
  PIN inner_wb_adr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END inner_wb_adr[14]
  PIN inner_wb_adr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END inner_wb_adr[15]
  PIN inner_wb_adr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END inner_wb_adr[16]
  PIN inner_wb_adr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END inner_wb_adr[17]
  PIN inner_wb_adr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END inner_wb_adr[18]
  PIN inner_wb_adr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END inner_wb_adr[19]
  PIN inner_wb_adr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END inner_wb_adr[1]
  PIN inner_wb_adr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END inner_wb_adr[20]
  PIN inner_wb_adr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END inner_wb_adr[21]
  PIN inner_wb_adr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END inner_wb_adr[22]
  PIN inner_wb_adr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END inner_wb_adr[23]
  PIN inner_wb_adr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END inner_wb_adr[2]
  PIN inner_wb_adr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END inner_wb_adr[3]
  PIN inner_wb_adr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END inner_wb_adr[4]
  PIN inner_wb_adr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END inner_wb_adr[5]
  PIN inner_wb_adr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END inner_wb_adr[6]
  PIN inner_wb_adr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END inner_wb_adr[7]
  PIN inner_wb_adr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END inner_wb_adr[8]
  PIN inner_wb_adr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END inner_wb_adr[9]
  PIN inner_wb_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END inner_wb_cyc
  PIN inner_wb_err
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END inner_wb_err
  PIN inner_wb_i_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END inner_wb_i_dat[0]
  PIN inner_wb_i_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END inner_wb_i_dat[10]
  PIN inner_wb_i_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END inner_wb_i_dat[11]
  PIN inner_wb_i_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END inner_wb_i_dat[12]
  PIN inner_wb_i_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END inner_wb_i_dat[13]
  PIN inner_wb_i_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END inner_wb_i_dat[14]
  PIN inner_wb_i_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END inner_wb_i_dat[15]
  PIN inner_wb_i_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END inner_wb_i_dat[1]
  PIN inner_wb_i_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END inner_wb_i_dat[2]
  PIN inner_wb_i_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END inner_wb_i_dat[3]
  PIN inner_wb_i_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END inner_wb_i_dat[4]
  PIN inner_wb_i_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END inner_wb_i_dat[5]
  PIN inner_wb_i_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END inner_wb_i_dat[6]
  PIN inner_wb_i_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END inner_wb_i_dat[7]
  PIN inner_wb_i_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END inner_wb_i_dat[8]
  PIN inner_wb_i_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END inner_wb_i_dat[9]
  PIN inner_wb_o_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END inner_wb_o_dat[0]
  PIN inner_wb_o_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END inner_wb_o_dat[10]
  PIN inner_wb_o_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END inner_wb_o_dat[11]
  PIN inner_wb_o_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END inner_wb_o_dat[12]
  PIN inner_wb_o_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END inner_wb_o_dat[13]
  PIN inner_wb_o_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END inner_wb_o_dat[14]
  PIN inner_wb_o_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END inner_wb_o_dat[15]
  PIN inner_wb_o_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END inner_wb_o_dat[1]
  PIN inner_wb_o_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END inner_wb_o_dat[2]
  PIN inner_wb_o_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END inner_wb_o_dat[3]
  PIN inner_wb_o_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END inner_wb_o_dat[4]
  PIN inner_wb_o_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END inner_wb_o_dat[5]
  PIN inner_wb_o_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END inner_wb_o_dat[6]
  PIN inner_wb_o_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END inner_wb_o_dat[7]
  PIN inner_wb_o_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END inner_wb_o_dat[8]
  PIN inner_wb_o_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END inner_wb_o_dat[9]
  PIN inner_wb_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END inner_wb_sel[0]
  PIN inner_wb_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END inner_wb_sel[1]
  PIN inner_wb_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END inner_wb_stb
  PIN inner_wb_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END inner_wb_we
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 788.885 ;
      LAYER met1 ;
        RECT 2.830 9.560 299.850 789.040 ;
      LAYER met2 ;
        RECT 2.860 4.280 299.820 788.985 ;
        RECT 2.860 4.000 6.710 4.280 ;
        RECT 7.550 4.000 10.850 4.280 ;
        RECT 11.690 4.000 14.990 4.280 ;
        RECT 15.830 4.000 19.130 4.280 ;
        RECT 19.970 4.000 23.270 4.280 ;
        RECT 24.110 4.000 27.410 4.280 ;
        RECT 28.250 4.000 31.550 4.280 ;
        RECT 32.390 4.000 35.690 4.280 ;
        RECT 36.530 4.000 39.830 4.280 ;
        RECT 40.670 4.000 43.970 4.280 ;
        RECT 44.810 4.000 48.110 4.280 ;
        RECT 48.950 4.000 52.250 4.280 ;
        RECT 53.090 4.000 56.390 4.280 ;
        RECT 57.230 4.000 60.530 4.280 ;
        RECT 61.370 4.000 64.670 4.280 ;
        RECT 65.510 4.000 68.810 4.280 ;
        RECT 69.650 4.000 72.950 4.280 ;
        RECT 73.790 4.000 77.090 4.280 ;
        RECT 77.930 4.000 81.230 4.280 ;
        RECT 82.070 4.000 85.370 4.280 ;
        RECT 86.210 4.000 89.510 4.280 ;
        RECT 90.350 4.000 93.650 4.280 ;
        RECT 94.490 4.000 97.790 4.280 ;
        RECT 98.630 4.000 101.930 4.280 ;
        RECT 102.770 4.000 106.070 4.280 ;
        RECT 106.910 4.000 110.210 4.280 ;
        RECT 111.050 4.000 114.350 4.280 ;
        RECT 115.190 4.000 118.490 4.280 ;
        RECT 119.330 4.000 122.630 4.280 ;
        RECT 123.470 4.000 126.770 4.280 ;
        RECT 127.610 4.000 130.910 4.280 ;
        RECT 131.750 4.000 135.050 4.280 ;
        RECT 135.890 4.000 139.190 4.280 ;
        RECT 140.030 4.000 143.330 4.280 ;
        RECT 144.170 4.000 147.470 4.280 ;
        RECT 148.310 4.000 151.610 4.280 ;
        RECT 152.450 4.000 155.750 4.280 ;
        RECT 156.590 4.000 159.890 4.280 ;
        RECT 160.730 4.000 164.030 4.280 ;
        RECT 164.870 4.000 168.170 4.280 ;
        RECT 169.010 4.000 172.310 4.280 ;
        RECT 173.150 4.000 176.450 4.280 ;
        RECT 177.290 4.000 180.590 4.280 ;
        RECT 181.430 4.000 184.730 4.280 ;
        RECT 185.570 4.000 188.870 4.280 ;
        RECT 189.710 4.000 193.010 4.280 ;
        RECT 193.850 4.000 197.150 4.280 ;
        RECT 197.990 4.000 201.290 4.280 ;
        RECT 202.130 4.000 205.430 4.280 ;
        RECT 206.270 4.000 209.570 4.280 ;
        RECT 210.410 4.000 213.710 4.280 ;
        RECT 214.550 4.000 217.850 4.280 ;
        RECT 218.690 4.000 221.990 4.280 ;
        RECT 222.830 4.000 226.130 4.280 ;
        RECT 226.970 4.000 230.270 4.280 ;
        RECT 231.110 4.000 234.410 4.280 ;
        RECT 235.250 4.000 238.550 4.280 ;
        RECT 239.390 4.000 242.690 4.280 ;
        RECT 243.530 4.000 246.830 4.280 ;
        RECT 247.670 4.000 250.970 4.280 ;
        RECT 251.810 4.000 255.110 4.280 ;
        RECT 255.950 4.000 259.250 4.280 ;
        RECT 260.090 4.000 263.390 4.280 ;
        RECT 264.230 4.000 267.530 4.280 ;
        RECT 268.370 4.000 271.670 4.280 ;
        RECT 272.510 4.000 275.810 4.280 ;
        RECT 276.650 4.000 279.950 4.280 ;
        RECT 280.790 4.000 284.090 4.280 ;
        RECT 284.930 4.000 288.230 4.280 ;
        RECT 289.070 4.000 292.370 4.280 ;
        RECT 293.210 4.000 299.820 4.280 ;
      LAYER met3 ;
        RECT 4.000 720.480 296.000 788.965 ;
        RECT 4.000 719.080 295.600 720.480 ;
        RECT 4.000 718.440 296.000 719.080 ;
        RECT 4.000 717.040 295.600 718.440 ;
        RECT 4.000 716.400 296.000 717.040 ;
        RECT 4.000 715.000 295.600 716.400 ;
        RECT 4.000 714.360 296.000 715.000 ;
        RECT 4.000 712.960 295.600 714.360 ;
        RECT 4.000 712.320 296.000 712.960 ;
        RECT 4.000 710.920 295.600 712.320 ;
        RECT 4.000 710.280 296.000 710.920 ;
        RECT 4.000 708.880 295.600 710.280 ;
        RECT 4.000 708.240 296.000 708.880 ;
        RECT 4.000 706.840 295.600 708.240 ;
        RECT 4.000 706.200 296.000 706.840 ;
        RECT 4.000 704.800 295.600 706.200 ;
        RECT 4.000 704.160 296.000 704.800 ;
        RECT 4.000 702.760 295.600 704.160 ;
        RECT 4.000 702.120 296.000 702.760 ;
        RECT 4.000 700.720 295.600 702.120 ;
        RECT 4.000 700.080 296.000 700.720 ;
        RECT 4.000 698.680 295.600 700.080 ;
        RECT 4.000 698.040 296.000 698.680 ;
        RECT 4.000 696.640 295.600 698.040 ;
        RECT 4.000 696.000 296.000 696.640 ;
        RECT 4.000 694.600 295.600 696.000 ;
        RECT 4.000 693.960 296.000 694.600 ;
        RECT 4.000 692.560 295.600 693.960 ;
        RECT 4.000 691.920 296.000 692.560 ;
        RECT 4.000 690.520 295.600 691.920 ;
        RECT 4.000 689.880 296.000 690.520 ;
        RECT 4.000 688.480 295.600 689.880 ;
        RECT 4.000 687.840 296.000 688.480 ;
        RECT 4.400 686.440 295.600 687.840 ;
        RECT 4.400 685.800 296.000 686.440 ;
        RECT 4.400 684.400 295.600 685.800 ;
        RECT 4.400 683.760 296.000 684.400 ;
        RECT 4.400 682.360 295.600 683.760 ;
        RECT 4.400 681.720 296.000 682.360 ;
        RECT 4.400 680.320 295.600 681.720 ;
        RECT 4.400 679.680 296.000 680.320 ;
        RECT 4.400 678.280 295.600 679.680 ;
        RECT 4.400 677.640 296.000 678.280 ;
        RECT 4.400 676.240 295.600 677.640 ;
        RECT 4.400 675.600 296.000 676.240 ;
        RECT 4.400 674.200 295.600 675.600 ;
        RECT 4.400 673.560 296.000 674.200 ;
        RECT 4.400 672.160 295.600 673.560 ;
        RECT 4.400 671.520 296.000 672.160 ;
        RECT 4.400 670.120 295.600 671.520 ;
        RECT 4.400 669.480 296.000 670.120 ;
        RECT 4.400 668.080 295.600 669.480 ;
        RECT 4.400 667.440 296.000 668.080 ;
        RECT 4.400 666.040 295.600 667.440 ;
        RECT 4.400 665.400 296.000 666.040 ;
        RECT 4.400 664.000 295.600 665.400 ;
        RECT 4.400 663.360 296.000 664.000 ;
        RECT 4.400 661.960 295.600 663.360 ;
        RECT 4.400 661.320 296.000 661.960 ;
        RECT 4.400 659.920 295.600 661.320 ;
        RECT 4.400 659.280 296.000 659.920 ;
        RECT 4.400 657.880 295.600 659.280 ;
        RECT 4.400 657.240 296.000 657.880 ;
        RECT 4.400 655.840 295.600 657.240 ;
        RECT 4.400 655.200 296.000 655.840 ;
        RECT 4.400 653.800 295.600 655.200 ;
        RECT 4.400 653.160 296.000 653.800 ;
        RECT 4.400 651.760 295.600 653.160 ;
        RECT 4.400 651.120 296.000 651.760 ;
        RECT 4.400 649.720 295.600 651.120 ;
        RECT 4.400 649.080 296.000 649.720 ;
        RECT 4.400 647.680 295.600 649.080 ;
        RECT 4.400 647.040 296.000 647.680 ;
        RECT 4.400 645.640 295.600 647.040 ;
        RECT 4.400 645.000 296.000 645.640 ;
        RECT 4.400 643.600 295.600 645.000 ;
        RECT 4.400 642.960 296.000 643.600 ;
        RECT 4.400 641.560 295.600 642.960 ;
        RECT 4.400 640.920 296.000 641.560 ;
        RECT 4.400 639.520 295.600 640.920 ;
        RECT 4.400 638.880 296.000 639.520 ;
        RECT 4.400 637.480 295.600 638.880 ;
        RECT 4.400 636.840 296.000 637.480 ;
        RECT 4.400 635.440 295.600 636.840 ;
        RECT 4.400 634.800 296.000 635.440 ;
        RECT 4.400 633.400 295.600 634.800 ;
        RECT 4.400 632.760 296.000 633.400 ;
        RECT 4.400 631.360 295.600 632.760 ;
        RECT 4.400 630.720 296.000 631.360 ;
        RECT 4.400 629.320 295.600 630.720 ;
        RECT 4.400 628.680 296.000 629.320 ;
        RECT 4.400 627.280 295.600 628.680 ;
        RECT 4.400 626.640 296.000 627.280 ;
        RECT 4.400 625.240 295.600 626.640 ;
        RECT 4.400 624.600 296.000 625.240 ;
        RECT 4.400 623.200 295.600 624.600 ;
        RECT 4.400 622.560 296.000 623.200 ;
        RECT 4.400 621.160 295.600 622.560 ;
        RECT 4.400 620.520 296.000 621.160 ;
        RECT 4.400 619.120 295.600 620.520 ;
        RECT 4.400 618.480 296.000 619.120 ;
        RECT 4.400 617.080 295.600 618.480 ;
        RECT 4.400 616.440 296.000 617.080 ;
        RECT 4.400 615.040 295.600 616.440 ;
        RECT 4.400 614.400 296.000 615.040 ;
        RECT 4.400 613.000 295.600 614.400 ;
        RECT 4.400 612.360 296.000 613.000 ;
        RECT 4.400 610.960 295.600 612.360 ;
        RECT 4.400 610.320 296.000 610.960 ;
        RECT 4.400 608.920 295.600 610.320 ;
        RECT 4.400 608.280 296.000 608.920 ;
        RECT 4.400 606.880 295.600 608.280 ;
        RECT 4.400 606.240 296.000 606.880 ;
        RECT 4.400 604.840 295.600 606.240 ;
        RECT 4.400 604.200 296.000 604.840 ;
        RECT 4.400 602.800 295.600 604.200 ;
        RECT 4.400 602.160 296.000 602.800 ;
        RECT 4.400 600.760 295.600 602.160 ;
        RECT 4.400 600.120 296.000 600.760 ;
        RECT 4.400 598.720 295.600 600.120 ;
        RECT 4.400 598.080 296.000 598.720 ;
        RECT 4.400 596.680 295.600 598.080 ;
        RECT 4.400 596.040 296.000 596.680 ;
        RECT 4.400 594.640 295.600 596.040 ;
        RECT 4.400 594.000 296.000 594.640 ;
        RECT 4.400 592.600 295.600 594.000 ;
        RECT 4.400 591.960 296.000 592.600 ;
        RECT 4.400 590.560 295.600 591.960 ;
        RECT 4.400 589.920 296.000 590.560 ;
        RECT 4.400 588.520 295.600 589.920 ;
        RECT 4.400 587.880 296.000 588.520 ;
        RECT 4.400 586.480 295.600 587.880 ;
        RECT 4.400 585.840 296.000 586.480 ;
        RECT 4.400 584.440 295.600 585.840 ;
        RECT 4.400 583.800 296.000 584.440 ;
        RECT 4.400 582.400 295.600 583.800 ;
        RECT 4.400 581.760 296.000 582.400 ;
        RECT 4.400 580.360 295.600 581.760 ;
        RECT 4.400 579.720 296.000 580.360 ;
        RECT 4.400 578.320 295.600 579.720 ;
        RECT 4.400 577.680 296.000 578.320 ;
        RECT 4.400 576.280 295.600 577.680 ;
        RECT 4.400 575.640 296.000 576.280 ;
        RECT 4.400 574.240 295.600 575.640 ;
        RECT 4.400 573.600 296.000 574.240 ;
        RECT 4.400 572.200 295.600 573.600 ;
        RECT 4.400 571.560 296.000 572.200 ;
        RECT 4.400 570.160 295.600 571.560 ;
        RECT 4.400 569.520 296.000 570.160 ;
        RECT 4.400 568.120 295.600 569.520 ;
        RECT 4.400 567.480 296.000 568.120 ;
        RECT 4.400 566.080 295.600 567.480 ;
        RECT 4.400 565.440 296.000 566.080 ;
        RECT 4.400 564.040 295.600 565.440 ;
        RECT 4.400 563.400 296.000 564.040 ;
        RECT 4.400 562.000 295.600 563.400 ;
        RECT 4.400 561.360 296.000 562.000 ;
        RECT 4.400 559.960 295.600 561.360 ;
        RECT 4.400 559.320 296.000 559.960 ;
        RECT 4.400 557.920 295.600 559.320 ;
        RECT 4.400 557.280 296.000 557.920 ;
        RECT 4.400 555.880 295.600 557.280 ;
        RECT 4.400 555.240 296.000 555.880 ;
        RECT 4.400 553.840 295.600 555.240 ;
        RECT 4.400 553.200 296.000 553.840 ;
        RECT 4.400 551.800 295.600 553.200 ;
        RECT 4.400 551.160 296.000 551.800 ;
        RECT 4.400 549.760 295.600 551.160 ;
        RECT 4.400 549.120 296.000 549.760 ;
        RECT 4.400 547.720 295.600 549.120 ;
        RECT 4.400 547.080 296.000 547.720 ;
        RECT 4.400 545.680 295.600 547.080 ;
        RECT 4.400 545.040 296.000 545.680 ;
        RECT 4.400 543.640 295.600 545.040 ;
        RECT 4.400 543.000 296.000 543.640 ;
        RECT 4.400 541.600 295.600 543.000 ;
        RECT 4.400 540.960 296.000 541.600 ;
        RECT 4.400 539.560 295.600 540.960 ;
        RECT 4.400 538.920 296.000 539.560 ;
        RECT 4.400 537.520 295.600 538.920 ;
        RECT 4.400 536.880 296.000 537.520 ;
        RECT 4.400 535.480 295.600 536.880 ;
        RECT 4.400 534.840 296.000 535.480 ;
        RECT 4.400 533.440 295.600 534.840 ;
        RECT 4.400 532.800 296.000 533.440 ;
        RECT 4.400 531.400 295.600 532.800 ;
        RECT 4.400 530.760 296.000 531.400 ;
        RECT 4.400 529.360 295.600 530.760 ;
        RECT 4.400 528.720 296.000 529.360 ;
        RECT 4.400 527.320 295.600 528.720 ;
        RECT 4.400 526.680 296.000 527.320 ;
        RECT 4.400 525.280 295.600 526.680 ;
        RECT 4.400 524.640 296.000 525.280 ;
        RECT 4.400 523.240 295.600 524.640 ;
        RECT 4.400 522.600 296.000 523.240 ;
        RECT 4.400 521.200 295.600 522.600 ;
        RECT 4.400 520.560 296.000 521.200 ;
        RECT 4.400 519.160 295.600 520.560 ;
        RECT 4.400 518.520 296.000 519.160 ;
        RECT 4.400 517.120 295.600 518.520 ;
        RECT 4.400 516.480 296.000 517.120 ;
        RECT 4.400 515.080 295.600 516.480 ;
        RECT 4.400 514.440 296.000 515.080 ;
        RECT 4.400 513.040 295.600 514.440 ;
        RECT 4.400 512.400 296.000 513.040 ;
        RECT 4.400 511.000 295.600 512.400 ;
        RECT 4.400 510.360 296.000 511.000 ;
        RECT 4.400 508.960 295.600 510.360 ;
        RECT 4.400 508.320 296.000 508.960 ;
        RECT 4.400 506.920 295.600 508.320 ;
        RECT 4.400 506.280 296.000 506.920 ;
        RECT 4.400 504.880 295.600 506.280 ;
        RECT 4.400 504.240 296.000 504.880 ;
        RECT 4.400 502.840 295.600 504.240 ;
        RECT 4.400 502.200 296.000 502.840 ;
        RECT 4.400 500.800 295.600 502.200 ;
        RECT 4.400 500.160 296.000 500.800 ;
        RECT 4.400 498.760 295.600 500.160 ;
        RECT 4.400 498.120 296.000 498.760 ;
        RECT 4.400 496.720 295.600 498.120 ;
        RECT 4.400 496.080 296.000 496.720 ;
        RECT 4.400 494.680 295.600 496.080 ;
        RECT 4.400 494.040 296.000 494.680 ;
        RECT 4.400 492.640 295.600 494.040 ;
        RECT 4.400 492.000 296.000 492.640 ;
        RECT 4.400 490.600 295.600 492.000 ;
        RECT 4.400 489.960 296.000 490.600 ;
        RECT 4.400 488.560 295.600 489.960 ;
        RECT 4.400 487.920 296.000 488.560 ;
        RECT 4.400 486.520 295.600 487.920 ;
        RECT 4.400 485.880 296.000 486.520 ;
        RECT 4.400 484.480 295.600 485.880 ;
        RECT 4.400 483.840 296.000 484.480 ;
        RECT 4.400 482.440 295.600 483.840 ;
        RECT 4.400 481.800 296.000 482.440 ;
        RECT 4.400 480.400 295.600 481.800 ;
        RECT 4.400 479.760 296.000 480.400 ;
        RECT 4.400 478.360 295.600 479.760 ;
        RECT 4.400 477.720 296.000 478.360 ;
        RECT 4.400 476.320 295.600 477.720 ;
        RECT 4.400 475.680 296.000 476.320 ;
        RECT 4.400 474.280 295.600 475.680 ;
        RECT 4.400 473.640 296.000 474.280 ;
        RECT 4.400 472.240 295.600 473.640 ;
        RECT 4.400 471.600 296.000 472.240 ;
        RECT 4.400 470.200 295.600 471.600 ;
        RECT 4.400 469.560 296.000 470.200 ;
        RECT 4.400 468.160 295.600 469.560 ;
        RECT 4.400 467.520 296.000 468.160 ;
        RECT 4.400 466.120 295.600 467.520 ;
        RECT 4.400 465.480 296.000 466.120 ;
        RECT 4.400 464.080 295.600 465.480 ;
        RECT 4.400 463.440 296.000 464.080 ;
        RECT 4.400 462.040 295.600 463.440 ;
        RECT 4.400 461.400 296.000 462.040 ;
        RECT 4.400 460.000 295.600 461.400 ;
        RECT 4.400 459.360 296.000 460.000 ;
        RECT 4.400 457.960 295.600 459.360 ;
        RECT 4.400 457.320 296.000 457.960 ;
        RECT 4.400 455.920 295.600 457.320 ;
        RECT 4.400 455.280 296.000 455.920 ;
        RECT 4.400 453.880 295.600 455.280 ;
        RECT 4.400 453.240 296.000 453.880 ;
        RECT 4.400 451.840 295.600 453.240 ;
        RECT 4.400 451.200 296.000 451.840 ;
        RECT 4.400 449.800 295.600 451.200 ;
        RECT 4.400 449.160 296.000 449.800 ;
        RECT 4.400 447.760 295.600 449.160 ;
        RECT 4.400 447.120 296.000 447.760 ;
        RECT 4.400 445.720 295.600 447.120 ;
        RECT 4.400 445.080 296.000 445.720 ;
        RECT 4.400 443.680 295.600 445.080 ;
        RECT 4.400 443.040 296.000 443.680 ;
        RECT 4.400 441.640 295.600 443.040 ;
        RECT 4.400 441.000 296.000 441.640 ;
        RECT 4.400 439.600 295.600 441.000 ;
        RECT 4.400 438.960 296.000 439.600 ;
        RECT 4.400 437.560 295.600 438.960 ;
        RECT 4.400 436.920 296.000 437.560 ;
        RECT 4.400 435.520 295.600 436.920 ;
        RECT 4.400 434.880 296.000 435.520 ;
        RECT 4.400 433.480 295.600 434.880 ;
        RECT 4.400 432.840 296.000 433.480 ;
        RECT 4.400 431.440 295.600 432.840 ;
        RECT 4.400 430.800 296.000 431.440 ;
        RECT 4.400 429.400 295.600 430.800 ;
        RECT 4.400 428.760 296.000 429.400 ;
        RECT 4.400 427.360 295.600 428.760 ;
        RECT 4.400 426.720 296.000 427.360 ;
        RECT 4.400 425.320 295.600 426.720 ;
        RECT 4.400 424.680 296.000 425.320 ;
        RECT 4.400 423.280 295.600 424.680 ;
        RECT 4.400 422.640 296.000 423.280 ;
        RECT 4.400 421.240 295.600 422.640 ;
        RECT 4.400 420.600 296.000 421.240 ;
        RECT 4.400 419.200 295.600 420.600 ;
        RECT 4.400 418.560 296.000 419.200 ;
        RECT 4.400 417.160 295.600 418.560 ;
        RECT 4.400 416.520 296.000 417.160 ;
        RECT 4.400 415.120 295.600 416.520 ;
        RECT 4.400 414.480 296.000 415.120 ;
        RECT 4.400 413.080 295.600 414.480 ;
        RECT 4.400 412.440 296.000 413.080 ;
        RECT 4.400 411.040 295.600 412.440 ;
        RECT 4.400 410.400 296.000 411.040 ;
        RECT 4.400 409.000 295.600 410.400 ;
        RECT 4.400 408.360 296.000 409.000 ;
        RECT 4.400 406.960 295.600 408.360 ;
        RECT 4.400 406.320 296.000 406.960 ;
        RECT 4.400 404.920 295.600 406.320 ;
        RECT 4.400 404.280 296.000 404.920 ;
        RECT 4.400 402.880 295.600 404.280 ;
        RECT 4.400 402.240 296.000 402.880 ;
        RECT 4.400 400.840 295.600 402.240 ;
        RECT 4.400 400.200 296.000 400.840 ;
        RECT 4.400 398.800 295.600 400.200 ;
        RECT 4.400 398.160 296.000 398.800 ;
        RECT 4.400 396.760 295.600 398.160 ;
        RECT 4.400 396.120 296.000 396.760 ;
        RECT 4.400 394.720 295.600 396.120 ;
        RECT 4.400 394.080 296.000 394.720 ;
        RECT 4.400 392.680 295.600 394.080 ;
        RECT 4.400 392.040 296.000 392.680 ;
        RECT 4.400 390.640 295.600 392.040 ;
        RECT 4.400 390.000 296.000 390.640 ;
        RECT 4.400 388.600 295.600 390.000 ;
        RECT 4.400 387.960 296.000 388.600 ;
        RECT 4.400 386.560 295.600 387.960 ;
        RECT 4.400 385.920 296.000 386.560 ;
        RECT 4.400 384.520 295.600 385.920 ;
        RECT 4.400 383.880 296.000 384.520 ;
        RECT 4.400 382.480 295.600 383.880 ;
        RECT 4.400 381.840 296.000 382.480 ;
        RECT 4.400 380.440 295.600 381.840 ;
        RECT 4.400 379.800 296.000 380.440 ;
        RECT 4.400 378.400 295.600 379.800 ;
        RECT 4.400 377.760 296.000 378.400 ;
        RECT 4.400 376.360 295.600 377.760 ;
        RECT 4.400 375.720 296.000 376.360 ;
        RECT 4.400 374.320 295.600 375.720 ;
        RECT 4.400 373.680 296.000 374.320 ;
        RECT 4.400 372.280 295.600 373.680 ;
        RECT 4.400 371.640 296.000 372.280 ;
        RECT 4.400 370.240 295.600 371.640 ;
        RECT 4.400 369.600 296.000 370.240 ;
        RECT 4.400 368.200 295.600 369.600 ;
        RECT 4.400 367.560 296.000 368.200 ;
        RECT 4.400 366.160 295.600 367.560 ;
        RECT 4.400 365.520 296.000 366.160 ;
        RECT 4.400 364.120 295.600 365.520 ;
        RECT 4.400 363.480 296.000 364.120 ;
        RECT 4.400 362.080 295.600 363.480 ;
        RECT 4.400 361.440 296.000 362.080 ;
        RECT 4.400 360.040 295.600 361.440 ;
        RECT 4.400 359.400 296.000 360.040 ;
        RECT 4.400 358.000 295.600 359.400 ;
        RECT 4.400 357.360 296.000 358.000 ;
        RECT 4.400 355.960 295.600 357.360 ;
        RECT 4.400 355.320 296.000 355.960 ;
        RECT 4.400 353.920 295.600 355.320 ;
        RECT 4.400 353.280 296.000 353.920 ;
        RECT 4.400 351.880 295.600 353.280 ;
        RECT 4.400 351.240 296.000 351.880 ;
        RECT 4.400 349.840 295.600 351.240 ;
        RECT 4.400 349.200 296.000 349.840 ;
        RECT 4.400 347.800 295.600 349.200 ;
        RECT 4.400 347.160 296.000 347.800 ;
        RECT 4.400 345.760 295.600 347.160 ;
        RECT 4.400 345.120 296.000 345.760 ;
        RECT 4.400 343.720 295.600 345.120 ;
        RECT 4.400 343.080 296.000 343.720 ;
        RECT 4.400 341.680 295.600 343.080 ;
        RECT 4.400 341.040 296.000 341.680 ;
        RECT 4.400 339.640 295.600 341.040 ;
        RECT 4.400 339.000 296.000 339.640 ;
        RECT 4.400 337.600 295.600 339.000 ;
        RECT 4.400 336.960 296.000 337.600 ;
        RECT 4.400 335.560 295.600 336.960 ;
        RECT 4.400 334.920 296.000 335.560 ;
        RECT 4.400 333.520 295.600 334.920 ;
        RECT 4.400 332.880 296.000 333.520 ;
        RECT 4.400 331.480 295.600 332.880 ;
        RECT 4.400 330.840 296.000 331.480 ;
        RECT 4.400 329.440 295.600 330.840 ;
        RECT 4.400 328.800 296.000 329.440 ;
        RECT 4.400 327.400 295.600 328.800 ;
        RECT 4.400 326.760 296.000 327.400 ;
        RECT 4.400 325.360 295.600 326.760 ;
        RECT 4.400 324.720 296.000 325.360 ;
        RECT 4.400 323.320 295.600 324.720 ;
        RECT 4.400 322.680 296.000 323.320 ;
        RECT 4.400 321.280 295.600 322.680 ;
        RECT 4.400 320.640 296.000 321.280 ;
        RECT 4.400 319.240 295.600 320.640 ;
        RECT 4.400 318.600 296.000 319.240 ;
        RECT 4.400 317.200 295.600 318.600 ;
        RECT 4.400 316.560 296.000 317.200 ;
        RECT 4.400 315.160 295.600 316.560 ;
        RECT 4.400 314.520 296.000 315.160 ;
        RECT 4.400 313.120 295.600 314.520 ;
        RECT 4.400 312.480 296.000 313.120 ;
        RECT 4.400 311.080 295.600 312.480 ;
        RECT 4.400 310.440 296.000 311.080 ;
        RECT 4.400 309.040 295.600 310.440 ;
        RECT 4.400 308.400 296.000 309.040 ;
        RECT 4.400 307.000 295.600 308.400 ;
        RECT 4.400 306.360 296.000 307.000 ;
        RECT 4.400 304.960 295.600 306.360 ;
        RECT 4.400 304.320 296.000 304.960 ;
        RECT 4.400 302.920 295.600 304.320 ;
        RECT 4.400 302.280 296.000 302.920 ;
        RECT 4.400 300.880 295.600 302.280 ;
        RECT 4.400 300.240 296.000 300.880 ;
        RECT 4.400 298.840 295.600 300.240 ;
        RECT 4.400 298.200 296.000 298.840 ;
        RECT 4.400 296.800 295.600 298.200 ;
        RECT 4.400 296.160 296.000 296.800 ;
        RECT 4.400 294.760 295.600 296.160 ;
        RECT 4.400 294.120 296.000 294.760 ;
        RECT 4.400 292.720 295.600 294.120 ;
        RECT 4.400 292.080 296.000 292.720 ;
        RECT 4.400 290.680 295.600 292.080 ;
        RECT 4.400 290.040 296.000 290.680 ;
        RECT 4.400 288.640 295.600 290.040 ;
        RECT 4.400 288.000 296.000 288.640 ;
        RECT 4.400 286.600 295.600 288.000 ;
        RECT 4.400 285.960 296.000 286.600 ;
        RECT 4.400 284.560 295.600 285.960 ;
        RECT 4.400 283.920 296.000 284.560 ;
        RECT 4.400 282.520 295.600 283.920 ;
        RECT 4.400 281.880 296.000 282.520 ;
        RECT 4.400 280.480 295.600 281.880 ;
        RECT 4.400 279.840 296.000 280.480 ;
        RECT 4.400 278.440 295.600 279.840 ;
        RECT 4.400 277.800 296.000 278.440 ;
        RECT 4.400 276.400 295.600 277.800 ;
        RECT 4.400 275.760 296.000 276.400 ;
        RECT 4.400 274.360 295.600 275.760 ;
        RECT 4.400 273.720 296.000 274.360 ;
        RECT 4.400 272.320 295.600 273.720 ;
        RECT 4.400 271.680 296.000 272.320 ;
        RECT 4.400 270.280 295.600 271.680 ;
        RECT 4.400 269.640 296.000 270.280 ;
        RECT 4.400 268.240 295.600 269.640 ;
        RECT 4.400 267.600 296.000 268.240 ;
        RECT 4.400 266.200 295.600 267.600 ;
        RECT 4.400 265.560 296.000 266.200 ;
        RECT 4.400 264.160 295.600 265.560 ;
        RECT 4.400 263.520 296.000 264.160 ;
        RECT 4.400 262.120 295.600 263.520 ;
        RECT 4.400 261.480 296.000 262.120 ;
        RECT 4.400 260.080 295.600 261.480 ;
        RECT 4.400 259.440 296.000 260.080 ;
        RECT 4.400 258.040 295.600 259.440 ;
        RECT 4.400 257.400 296.000 258.040 ;
        RECT 4.400 256.000 295.600 257.400 ;
        RECT 4.400 255.360 296.000 256.000 ;
        RECT 4.400 253.960 295.600 255.360 ;
        RECT 4.400 253.320 296.000 253.960 ;
        RECT 4.400 251.920 295.600 253.320 ;
        RECT 4.400 251.280 296.000 251.920 ;
        RECT 4.400 249.880 295.600 251.280 ;
        RECT 4.400 249.240 296.000 249.880 ;
        RECT 4.400 247.840 295.600 249.240 ;
        RECT 4.400 247.200 296.000 247.840 ;
        RECT 4.400 245.800 295.600 247.200 ;
        RECT 4.400 245.160 296.000 245.800 ;
        RECT 4.400 243.760 295.600 245.160 ;
        RECT 4.400 243.120 296.000 243.760 ;
        RECT 4.400 241.720 295.600 243.120 ;
        RECT 4.400 241.080 296.000 241.720 ;
        RECT 4.400 239.680 295.600 241.080 ;
        RECT 4.400 239.040 296.000 239.680 ;
        RECT 4.400 237.640 295.600 239.040 ;
        RECT 4.400 237.000 296.000 237.640 ;
        RECT 4.400 235.600 295.600 237.000 ;
        RECT 4.400 234.960 296.000 235.600 ;
        RECT 4.400 233.560 295.600 234.960 ;
        RECT 4.400 232.920 296.000 233.560 ;
        RECT 4.400 231.520 295.600 232.920 ;
        RECT 4.400 230.880 296.000 231.520 ;
        RECT 4.400 229.480 295.600 230.880 ;
        RECT 4.400 228.840 296.000 229.480 ;
        RECT 4.400 227.440 295.600 228.840 ;
        RECT 4.400 226.800 296.000 227.440 ;
        RECT 4.400 225.400 295.600 226.800 ;
        RECT 4.400 224.760 296.000 225.400 ;
        RECT 4.400 223.360 295.600 224.760 ;
        RECT 4.400 222.720 296.000 223.360 ;
        RECT 4.400 221.320 295.600 222.720 ;
        RECT 4.400 220.680 296.000 221.320 ;
        RECT 4.400 219.280 295.600 220.680 ;
        RECT 4.400 218.640 296.000 219.280 ;
        RECT 4.400 217.240 295.600 218.640 ;
        RECT 4.400 216.600 296.000 217.240 ;
        RECT 4.400 215.200 295.600 216.600 ;
        RECT 4.400 214.560 296.000 215.200 ;
        RECT 4.400 213.160 295.600 214.560 ;
        RECT 4.400 212.520 296.000 213.160 ;
        RECT 4.400 211.120 295.600 212.520 ;
        RECT 4.400 210.480 296.000 211.120 ;
        RECT 4.400 209.080 295.600 210.480 ;
        RECT 4.400 208.440 296.000 209.080 ;
        RECT 4.400 207.040 295.600 208.440 ;
        RECT 4.400 206.400 296.000 207.040 ;
        RECT 4.400 205.000 295.600 206.400 ;
        RECT 4.400 204.360 296.000 205.000 ;
        RECT 4.400 202.960 295.600 204.360 ;
        RECT 4.400 202.320 296.000 202.960 ;
        RECT 4.400 200.920 295.600 202.320 ;
        RECT 4.400 200.280 296.000 200.920 ;
        RECT 4.400 198.880 295.600 200.280 ;
        RECT 4.400 198.240 296.000 198.880 ;
        RECT 4.400 196.840 295.600 198.240 ;
        RECT 4.400 196.200 296.000 196.840 ;
        RECT 4.400 194.800 295.600 196.200 ;
        RECT 4.400 194.160 296.000 194.800 ;
        RECT 4.400 192.760 295.600 194.160 ;
        RECT 4.400 192.120 296.000 192.760 ;
        RECT 4.400 190.720 295.600 192.120 ;
        RECT 4.400 190.080 296.000 190.720 ;
        RECT 4.400 188.680 295.600 190.080 ;
        RECT 4.400 188.040 296.000 188.680 ;
        RECT 4.400 186.640 295.600 188.040 ;
        RECT 4.400 186.000 296.000 186.640 ;
        RECT 4.400 184.600 295.600 186.000 ;
        RECT 4.400 183.960 296.000 184.600 ;
        RECT 4.400 182.560 295.600 183.960 ;
        RECT 4.400 181.920 296.000 182.560 ;
        RECT 4.400 180.520 295.600 181.920 ;
        RECT 4.400 179.880 296.000 180.520 ;
        RECT 4.400 178.480 295.600 179.880 ;
        RECT 4.400 177.840 296.000 178.480 ;
        RECT 4.400 176.440 295.600 177.840 ;
        RECT 4.400 175.800 296.000 176.440 ;
        RECT 4.400 174.400 295.600 175.800 ;
        RECT 4.400 173.760 296.000 174.400 ;
        RECT 4.400 172.360 295.600 173.760 ;
        RECT 4.400 171.720 296.000 172.360 ;
        RECT 4.400 170.320 295.600 171.720 ;
        RECT 4.400 169.680 296.000 170.320 ;
        RECT 4.400 168.280 295.600 169.680 ;
        RECT 4.400 167.640 296.000 168.280 ;
        RECT 4.400 166.240 295.600 167.640 ;
        RECT 4.400 165.600 296.000 166.240 ;
        RECT 4.400 164.200 295.600 165.600 ;
        RECT 4.400 163.560 296.000 164.200 ;
        RECT 4.400 162.160 295.600 163.560 ;
        RECT 4.400 161.520 296.000 162.160 ;
        RECT 4.400 160.120 295.600 161.520 ;
        RECT 4.400 159.480 296.000 160.120 ;
        RECT 4.400 158.080 295.600 159.480 ;
        RECT 4.400 157.440 296.000 158.080 ;
        RECT 4.400 156.040 295.600 157.440 ;
        RECT 4.400 155.400 296.000 156.040 ;
        RECT 4.400 154.000 295.600 155.400 ;
        RECT 4.400 153.360 296.000 154.000 ;
        RECT 4.400 151.960 295.600 153.360 ;
        RECT 4.400 151.320 296.000 151.960 ;
        RECT 4.400 149.920 295.600 151.320 ;
        RECT 4.400 149.280 296.000 149.920 ;
        RECT 4.400 147.880 295.600 149.280 ;
        RECT 4.400 147.240 296.000 147.880 ;
        RECT 4.400 145.840 295.600 147.240 ;
        RECT 4.400 145.200 296.000 145.840 ;
        RECT 4.400 143.800 295.600 145.200 ;
        RECT 4.400 143.160 296.000 143.800 ;
        RECT 4.400 141.760 295.600 143.160 ;
        RECT 4.400 141.120 296.000 141.760 ;
        RECT 4.400 139.720 295.600 141.120 ;
        RECT 4.400 139.080 296.000 139.720 ;
        RECT 4.400 137.680 295.600 139.080 ;
        RECT 4.400 137.040 296.000 137.680 ;
        RECT 4.400 135.640 295.600 137.040 ;
        RECT 4.400 135.000 296.000 135.640 ;
        RECT 4.400 133.600 295.600 135.000 ;
        RECT 4.400 132.960 296.000 133.600 ;
        RECT 4.400 131.560 295.600 132.960 ;
        RECT 4.400 130.920 296.000 131.560 ;
        RECT 4.400 129.520 295.600 130.920 ;
        RECT 4.400 128.880 296.000 129.520 ;
        RECT 4.400 127.480 295.600 128.880 ;
        RECT 4.400 126.840 296.000 127.480 ;
        RECT 4.400 125.440 295.600 126.840 ;
        RECT 4.400 124.800 296.000 125.440 ;
        RECT 4.400 123.400 295.600 124.800 ;
        RECT 4.400 122.760 296.000 123.400 ;
        RECT 4.400 121.360 295.600 122.760 ;
        RECT 4.400 120.720 296.000 121.360 ;
        RECT 4.400 119.320 295.600 120.720 ;
        RECT 4.400 118.680 296.000 119.320 ;
        RECT 4.400 117.280 295.600 118.680 ;
        RECT 4.400 116.640 296.000 117.280 ;
        RECT 4.400 115.240 295.600 116.640 ;
        RECT 4.400 114.600 296.000 115.240 ;
        RECT 4.400 113.200 295.600 114.600 ;
        RECT 4.400 112.560 296.000 113.200 ;
        RECT 4.400 111.160 295.600 112.560 ;
        RECT 4.000 110.520 296.000 111.160 ;
        RECT 4.000 109.120 295.600 110.520 ;
        RECT 4.000 108.480 296.000 109.120 ;
        RECT 4.000 107.080 295.600 108.480 ;
        RECT 4.000 106.440 296.000 107.080 ;
        RECT 4.000 105.040 295.600 106.440 ;
        RECT 4.000 104.400 296.000 105.040 ;
        RECT 4.000 103.000 295.600 104.400 ;
        RECT 4.000 102.360 296.000 103.000 ;
        RECT 4.000 100.960 295.600 102.360 ;
        RECT 4.000 100.320 296.000 100.960 ;
        RECT 4.000 98.920 295.600 100.320 ;
        RECT 4.000 98.280 296.000 98.920 ;
        RECT 4.000 96.880 295.600 98.280 ;
        RECT 4.000 96.240 296.000 96.880 ;
        RECT 4.000 94.840 295.600 96.240 ;
        RECT 4.000 94.200 296.000 94.840 ;
        RECT 4.000 92.800 295.600 94.200 ;
        RECT 4.000 92.160 296.000 92.800 ;
        RECT 4.000 90.760 295.600 92.160 ;
        RECT 4.000 90.120 296.000 90.760 ;
        RECT 4.000 88.720 295.600 90.120 ;
        RECT 4.000 88.080 296.000 88.720 ;
        RECT 4.000 86.680 295.600 88.080 ;
        RECT 4.000 86.040 296.000 86.680 ;
        RECT 4.000 84.640 295.600 86.040 ;
        RECT 4.000 84.000 296.000 84.640 ;
        RECT 4.000 82.600 295.600 84.000 ;
        RECT 4.000 81.960 296.000 82.600 ;
        RECT 4.000 80.560 295.600 81.960 ;
        RECT 4.000 79.920 296.000 80.560 ;
        RECT 4.000 78.520 295.600 79.920 ;
        RECT 4.000 10.715 296.000 78.520 ;
      LAYER met4 ;
        RECT 2.150 11.735 20.640 757.345 ;
        RECT 23.040 11.735 97.440 757.345 ;
        RECT 99.840 11.735 174.240 757.345 ;
        RECT 176.640 11.735 251.040 757.345 ;
        RECT 253.440 11.735 288.585 757.345 ;
  END
END interconnect_inner
END LIBRARY

