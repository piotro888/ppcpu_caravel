magic
tech sky130B
magscale 1 2
timestamp 1663070243
<< obsli1 >>
rect 1104 2159 38824 47345
<< obsm1 >>
rect 14 1708 39362 47524
<< metal2 >>
rect 18 49200 74 50000
rect 662 49200 718 50000
rect 1306 49200 1362 50000
rect 1950 49200 2006 50000
rect 2594 49200 2650 50000
rect 3238 49200 3294 50000
rect 3882 49200 3938 50000
rect 4526 49200 4582 50000
rect 5170 49200 5226 50000
rect 5814 49200 5870 50000
rect 6458 49200 6514 50000
rect 7102 49200 7158 50000
rect 7746 49200 7802 50000
rect 8390 49200 8446 50000
rect 9034 49200 9090 50000
rect 9678 49200 9734 50000
rect 10966 49200 11022 50000
rect 11610 49200 11666 50000
rect 12254 49200 12310 50000
rect 12898 49200 12954 50000
rect 13542 49200 13598 50000
rect 14186 49200 14242 50000
rect 14830 49200 14886 50000
rect 15474 49200 15530 50000
rect 16118 49200 16174 50000
rect 16762 49200 16818 50000
rect 17406 49200 17462 50000
rect 18050 49200 18106 50000
rect 18694 49200 18750 50000
rect 19338 49200 19394 50000
rect 19982 49200 20038 50000
rect 20626 49200 20682 50000
rect 21270 49200 21326 50000
rect 21914 49200 21970 50000
rect 22558 49200 22614 50000
rect 23202 49200 23258 50000
rect 23846 49200 23902 50000
rect 24490 49200 24546 50000
rect 25778 49200 25834 50000
rect 26422 49200 26478 50000
rect 27066 49200 27122 50000
rect 27710 49200 27766 50000
rect 28354 49200 28410 50000
rect 28998 49200 29054 50000
rect 29642 49200 29698 50000
rect 30286 49200 30342 50000
rect 30930 49200 30986 50000
rect 31574 49200 31630 50000
rect 32218 49200 32274 50000
rect 32862 49200 32918 50000
rect 33506 49200 33562 50000
rect 34150 49200 34206 50000
rect 34794 49200 34850 50000
rect 35438 49200 35494 50000
rect 36082 49200 36138 50000
rect 36726 49200 36782 50000
rect 37370 49200 37426 50000
rect 38014 49200 38070 50000
rect 38658 49200 38714 50000
rect 39302 49200 39358 50000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
<< obsm2 >>
rect 130 49144 606 49745
rect 774 49144 1250 49745
rect 1418 49144 1894 49745
rect 2062 49144 2538 49745
rect 2706 49144 3182 49745
rect 3350 49144 3826 49745
rect 3994 49144 4470 49745
rect 4638 49144 5114 49745
rect 5282 49144 5758 49745
rect 5926 49144 6402 49745
rect 6570 49144 7046 49745
rect 7214 49144 7690 49745
rect 7858 49144 8334 49745
rect 8502 49144 8978 49745
rect 9146 49144 9622 49745
rect 9790 49144 10910 49745
rect 11078 49144 11554 49745
rect 11722 49144 12198 49745
rect 12366 49144 12842 49745
rect 13010 49144 13486 49745
rect 13654 49144 14130 49745
rect 14298 49144 14774 49745
rect 14942 49144 15418 49745
rect 15586 49144 16062 49745
rect 16230 49144 16706 49745
rect 16874 49144 17350 49745
rect 17518 49144 17994 49745
rect 18162 49144 18638 49745
rect 18806 49144 19282 49745
rect 19450 49144 19926 49745
rect 20094 49144 20570 49745
rect 20738 49144 21214 49745
rect 21382 49144 21858 49745
rect 22026 49144 22502 49745
rect 22670 49144 23146 49745
rect 23314 49144 23790 49745
rect 23958 49144 24434 49745
rect 24602 49144 25722 49745
rect 25890 49144 26366 49745
rect 26534 49144 27010 49745
rect 27178 49144 27654 49745
rect 27822 49144 28298 49745
rect 28466 49144 28942 49745
rect 29110 49144 29586 49745
rect 29754 49144 30230 49745
rect 30398 49144 30874 49745
rect 31042 49144 31518 49745
rect 31686 49144 32162 49745
rect 32330 49144 32806 49745
rect 32974 49144 33450 49745
rect 33618 49144 34094 49745
rect 34262 49144 34738 49745
rect 34906 49144 35382 49745
rect 35550 49144 36026 49745
rect 36194 49144 36670 49745
rect 36838 49144 37314 49745
rect 37482 49144 37958 49745
rect 38126 49144 38602 49745
rect 38770 49144 39246 49745
rect 20 856 39356 49144
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 1894 856
rect 2062 31 2538 856
rect 2706 31 3182 856
rect 3350 31 3826 856
rect 3994 31 4470 856
rect 4638 31 5114 856
rect 5282 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7046 856
rect 7214 31 7690 856
rect 7858 31 8334 856
rect 8502 31 8978 856
rect 9146 31 9622 856
rect 9790 31 10266 856
rect 10434 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12198 856
rect 12366 31 12842 856
rect 13010 31 13486 856
rect 13654 31 14774 856
rect 14942 31 15418 856
rect 15586 31 16062 856
rect 16230 31 16706 856
rect 16874 31 17350 856
rect 17518 31 17994 856
rect 18162 31 18638 856
rect 18806 31 19282 856
rect 19450 31 19926 856
rect 20094 31 20570 856
rect 20738 31 21214 856
rect 21382 31 21858 856
rect 22026 31 22502 856
rect 22670 31 23146 856
rect 23314 31 23790 856
rect 23958 31 24434 856
rect 24602 31 25078 856
rect 25246 31 25722 856
rect 25890 31 26366 856
rect 26534 31 27010 856
rect 27178 31 27654 856
rect 27822 31 28298 856
rect 28466 31 29586 856
rect 29754 31 30230 856
rect 30398 31 30874 856
rect 31042 31 31518 856
rect 31686 31 32162 856
rect 32330 31 32806 856
rect 32974 31 33450 856
rect 33618 31 34094 856
rect 34262 31 34738 856
rect 34906 31 35382 856
rect 35550 31 36026 856
rect 36194 31 36670 856
rect 36838 31 37314 856
rect 37482 31 37958 856
rect 38126 31 38602 856
rect 38770 31 39246 856
<< metal3 >>
rect 0 49648 800 49768
rect 0 48968 800 49088
rect 39200 48968 40000 49088
rect 0 48288 800 48408
rect 39200 48288 40000 48408
rect 0 47608 800 47728
rect 39200 47608 40000 47728
rect 0 46928 800 47048
rect 39200 46928 40000 47048
rect 39200 46248 40000 46368
rect 0 45568 800 45688
rect 39200 45568 40000 45688
rect 0 44888 800 45008
rect 39200 44888 40000 45008
rect 0 44208 800 44328
rect 39200 44208 40000 44328
rect 0 43528 800 43648
rect 39200 43528 40000 43648
rect 0 42848 800 42968
rect 39200 42848 40000 42968
rect 0 42168 800 42288
rect 39200 42168 40000 42288
rect 0 41488 800 41608
rect 39200 41488 40000 41608
rect 0 40808 800 40928
rect 39200 40808 40000 40928
rect 0 40128 800 40248
rect 39200 40128 40000 40248
rect 0 39448 800 39568
rect 39200 39448 40000 39568
rect 0 38768 800 38888
rect 39200 38768 40000 38888
rect 0 38088 800 38208
rect 39200 38088 40000 38208
rect 0 37408 800 37528
rect 39200 37408 40000 37528
rect 0 36728 800 36848
rect 39200 36728 40000 36848
rect 0 36048 800 36168
rect 39200 36048 40000 36168
rect 0 35368 800 35488
rect 39200 35368 40000 35488
rect 0 34688 800 34808
rect 0 34008 800 34128
rect 39200 34008 40000 34128
rect 0 33328 800 33448
rect 39200 33328 40000 33448
rect 0 32648 800 32768
rect 39200 32648 40000 32768
rect 0 31968 800 32088
rect 39200 31968 40000 32088
rect 0 31288 800 31408
rect 39200 31288 40000 31408
rect 39200 30608 40000 30728
rect 0 29928 800 30048
rect 39200 29928 40000 30048
rect 0 29248 800 29368
rect 39200 29248 40000 29368
rect 0 28568 800 28688
rect 39200 28568 40000 28688
rect 0 27888 800 28008
rect 39200 27888 40000 28008
rect 0 27208 800 27328
rect 39200 27208 40000 27328
rect 0 26528 800 26648
rect 39200 26528 40000 26648
rect 0 25848 800 25968
rect 39200 25848 40000 25968
rect 0 25168 800 25288
rect 39200 25168 40000 25288
rect 0 24488 800 24608
rect 39200 24488 40000 24608
rect 0 23808 800 23928
rect 39200 23808 40000 23928
rect 0 23128 800 23248
rect 39200 23128 40000 23248
rect 0 22448 800 22568
rect 39200 22448 40000 22568
rect 0 21768 800 21888
rect 39200 21768 40000 21888
rect 0 21088 800 21208
rect 39200 21088 40000 21208
rect 0 20408 800 20528
rect 39200 20408 40000 20528
rect 0 19728 800 19848
rect 39200 19728 40000 19848
rect 0 19048 800 19168
rect 0 18368 800 18488
rect 39200 18368 40000 18488
rect 0 17688 800 17808
rect 39200 17688 40000 17808
rect 0 17008 800 17128
rect 39200 17008 40000 17128
rect 0 16328 800 16448
rect 39200 16328 40000 16448
rect 0 15648 800 15768
rect 39200 15648 40000 15768
rect 39200 14968 40000 15088
rect 0 14288 800 14408
rect 39200 14288 40000 14408
rect 0 13608 800 13728
rect 39200 13608 40000 13728
rect 0 12928 800 13048
rect 39200 12928 40000 13048
rect 0 12248 800 12368
rect 39200 12248 40000 12368
rect 0 11568 800 11688
rect 39200 11568 40000 11688
rect 0 10888 800 11008
rect 39200 10888 40000 11008
rect 0 10208 800 10328
rect 39200 10208 40000 10328
rect 0 9528 800 9648
rect 39200 9528 40000 9648
rect 0 8848 800 8968
rect 39200 8848 40000 8968
rect 0 8168 800 8288
rect 39200 8168 40000 8288
rect 0 7488 800 7608
rect 39200 7488 40000 7608
rect 0 6808 800 6928
rect 39200 6808 40000 6928
rect 0 6128 800 6248
rect 39200 6128 40000 6248
rect 0 5448 800 5568
rect 39200 5448 40000 5568
rect 0 4768 800 4888
rect 39200 4768 40000 4888
rect 0 4088 800 4208
rect 39200 4088 40000 4208
rect 0 3408 800 3528
rect 0 2728 800 2848
rect 39200 2728 40000 2848
rect 0 2048 800 2168
rect 39200 2048 40000 2168
rect 0 1368 800 1488
rect 39200 1368 40000 1488
rect 0 688 800 808
rect 39200 688 40000 808
rect 39200 8 40000 128
<< obsm3 >>
rect 880 49568 39200 49741
rect 800 49168 39200 49568
rect 880 48888 39120 49168
rect 800 48488 39200 48888
rect 880 48208 39120 48488
rect 800 47808 39200 48208
rect 880 47528 39120 47808
rect 800 47128 39200 47528
rect 880 46848 39120 47128
rect 800 46448 39200 46848
rect 800 46168 39120 46448
rect 800 45768 39200 46168
rect 880 45488 39120 45768
rect 800 45088 39200 45488
rect 880 44808 39120 45088
rect 800 44408 39200 44808
rect 880 44128 39120 44408
rect 800 43728 39200 44128
rect 880 43448 39120 43728
rect 800 43048 39200 43448
rect 880 42768 39120 43048
rect 800 42368 39200 42768
rect 880 42088 39120 42368
rect 800 41688 39200 42088
rect 880 41408 39120 41688
rect 800 41008 39200 41408
rect 880 40728 39120 41008
rect 800 40328 39200 40728
rect 880 40048 39120 40328
rect 800 39648 39200 40048
rect 880 39368 39120 39648
rect 800 38968 39200 39368
rect 880 38688 39120 38968
rect 800 38288 39200 38688
rect 880 38008 39120 38288
rect 800 37608 39200 38008
rect 880 37328 39120 37608
rect 800 36928 39200 37328
rect 880 36648 39120 36928
rect 800 36248 39200 36648
rect 880 35968 39120 36248
rect 800 35568 39200 35968
rect 880 35288 39120 35568
rect 800 34888 39200 35288
rect 880 34608 39200 34888
rect 800 34208 39200 34608
rect 880 33928 39120 34208
rect 800 33528 39200 33928
rect 880 33248 39120 33528
rect 800 32848 39200 33248
rect 880 32568 39120 32848
rect 800 32168 39200 32568
rect 880 31888 39120 32168
rect 800 31488 39200 31888
rect 880 31208 39120 31488
rect 800 30808 39200 31208
rect 800 30528 39120 30808
rect 800 30128 39200 30528
rect 880 29848 39120 30128
rect 800 29448 39200 29848
rect 880 29168 39120 29448
rect 800 28768 39200 29168
rect 880 28488 39120 28768
rect 800 28088 39200 28488
rect 880 27808 39120 28088
rect 800 27408 39200 27808
rect 880 27128 39120 27408
rect 800 26728 39200 27128
rect 880 26448 39120 26728
rect 800 26048 39200 26448
rect 880 25768 39120 26048
rect 800 25368 39200 25768
rect 880 25088 39120 25368
rect 800 24688 39200 25088
rect 880 24408 39120 24688
rect 800 24008 39200 24408
rect 880 23728 39120 24008
rect 800 23328 39200 23728
rect 880 23048 39120 23328
rect 800 22648 39200 23048
rect 880 22368 39120 22648
rect 800 21968 39200 22368
rect 880 21688 39120 21968
rect 800 21288 39200 21688
rect 880 21008 39120 21288
rect 800 20608 39200 21008
rect 880 20328 39120 20608
rect 800 19928 39200 20328
rect 880 19648 39120 19928
rect 800 19248 39200 19648
rect 880 18968 39200 19248
rect 800 18568 39200 18968
rect 880 18288 39120 18568
rect 800 17888 39200 18288
rect 880 17608 39120 17888
rect 800 17208 39200 17608
rect 880 16928 39120 17208
rect 800 16528 39200 16928
rect 880 16248 39120 16528
rect 800 15848 39200 16248
rect 880 15568 39120 15848
rect 800 15168 39200 15568
rect 800 14888 39120 15168
rect 800 14488 39200 14888
rect 880 14208 39120 14488
rect 800 13808 39200 14208
rect 880 13528 39120 13808
rect 800 13128 39200 13528
rect 880 12848 39120 13128
rect 800 12448 39200 12848
rect 880 12168 39120 12448
rect 800 11768 39200 12168
rect 880 11488 39120 11768
rect 800 11088 39200 11488
rect 880 10808 39120 11088
rect 800 10408 39200 10808
rect 880 10128 39120 10408
rect 800 9728 39200 10128
rect 880 9448 39120 9728
rect 800 9048 39200 9448
rect 880 8768 39120 9048
rect 800 8368 39200 8768
rect 880 8088 39120 8368
rect 800 7688 39200 8088
rect 880 7408 39120 7688
rect 800 7008 39200 7408
rect 880 6728 39120 7008
rect 800 6328 39200 6728
rect 880 6048 39120 6328
rect 800 5648 39200 6048
rect 880 5368 39120 5648
rect 800 4968 39200 5368
rect 880 4688 39120 4968
rect 800 4288 39200 4688
rect 880 4008 39120 4288
rect 800 3608 39200 4008
rect 880 3328 39200 3608
rect 800 2928 39200 3328
rect 880 2648 39120 2928
rect 800 2248 39200 2648
rect 880 1968 39120 2248
rect 800 1568 39200 1968
rect 880 1288 39120 1568
rect 800 888 39200 1288
rect 880 608 39120 888
rect 800 208 39200 608
rect 800 35 39120 208
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
<< labels >>
rlabel metal3 s 0 47608 800 47728 6 c_wb_4_burst
port 1 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 c_wb_8_burst
port 2 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 c_wb_ack_cmp
port 3 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 c_wb_adr[0]
port 4 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 c_wb_adr[10]
port 5 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 c_wb_adr[11]
port 6 nsew signal output
rlabel metal3 s 39200 27208 40000 27328 6 c_wb_adr[12]
port 7 nsew signal output
rlabel metal2 s 15474 49200 15530 50000 6 c_wb_adr[13]
port 8 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 c_wb_adr[14]
port 9 nsew signal output
rlabel metal3 s 39200 15648 40000 15768 6 c_wb_adr[15]
port 10 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 c_wb_adr[16]
port 11 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 c_wb_adr[17]
port 12 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 c_wb_adr[18]
port 13 nsew signal output
rlabel metal2 s 7746 49200 7802 50000 6 c_wb_adr[19]
port 14 nsew signal output
rlabel metal3 s 39200 36048 40000 36168 6 c_wb_adr[1]
port 15 nsew signal output
rlabel metal2 s 27710 49200 27766 50000 6 c_wb_adr[20]
port 16 nsew signal output
rlabel metal3 s 39200 29928 40000 30048 6 c_wb_adr[21]
port 17 nsew signal output
rlabel metal3 s 39200 27888 40000 28008 6 c_wb_adr[22]
port 18 nsew signal output
rlabel metal3 s 39200 6128 40000 6248 6 c_wb_adr[23]
port 19 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 c_wb_adr[2]
port 20 nsew signal output
rlabel metal2 s 27066 49200 27122 50000 6 c_wb_adr[3]
port 21 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 c_wb_adr[4]
port 22 nsew signal output
rlabel metal2 s 26422 49200 26478 50000 6 c_wb_adr[5]
port 23 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 c_wb_adr[6]
port 24 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 c_wb_adr[7]
port 25 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 c_wb_adr[8]
port 26 nsew signal output
rlabel metal3 s 39200 23808 40000 23928 6 c_wb_adr[9]
port 27 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 c_wb_cyc
port 28 nsew signal output
rlabel metal2 s 8390 49200 8446 50000 6 c_wb_err_cmp
port 29 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 c_wb_i_dat_cmp[0]
port 30 nsew signal input
rlabel metal2 s 35438 49200 35494 50000 6 c_wb_i_dat_cmp[10]
port 31 nsew signal input
rlabel metal3 s 39200 45568 40000 45688 6 c_wb_i_dat_cmp[11]
port 32 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 c_wb_i_dat_cmp[12]
port 33 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 c_wb_i_dat_cmp[13]
port 34 nsew signal input
rlabel metal2 s 6458 49200 6514 50000 6 c_wb_i_dat_cmp[14]
port 35 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 c_wb_i_dat_cmp[15]
port 36 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 c_wb_i_dat_cmp[1]
port 37 nsew signal input
rlabel metal3 s 39200 31288 40000 31408 6 c_wb_i_dat_cmp[2]
port 38 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 c_wb_i_dat_cmp[3]
port 39 nsew signal input
rlabel metal2 s 3882 49200 3938 50000 6 c_wb_i_dat_cmp[4]
port 40 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 c_wb_i_dat_cmp[5]
port 41 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 c_wb_i_dat_cmp[6]
port 42 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 c_wb_i_dat_cmp[7]
port 43 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 c_wb_i_dat_cmp[8]
port 44 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 c_wb_i_dat_cmp[9]
port 45 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 c_wb_o_dat[0]
port 46 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 c_wb_o_dat[10]
port 47 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 c_wb_o_dat[11]
port 48 nsew signal output
rlabel metal2 s 17406 49200 17462 50000 6 c_wb_o_dat[12]
port 49 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 c_wb_o_dat[13]
port 50 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 c_wb_o_dat[14]
port 51 nsew signal output
rlabel metal3 s 39200 4768 40000 4888 6 c_wb_o_dat[15]
port 52 nsew signal output
rlabel metal2 s 30286 49200 30342 50000 6 c_wb_o_dat[1]
port 53 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 c_wb_o_dat[2]
port 54 nsew signal output
rlabel metal2 s 9678 49200 9734 50000 6 c_wb_o_dat[3]
port 55 nsew signal output
rlabel metal2 s 662 49200 718 50000 6 c_wb_o_dat[4]
port 56 nsew signal output
rlabel metal3 s 39200 1368 40000 1488 6 c_wb_o_dat[5]
port 57 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 c_wb_o_dat[6]
port 58 nsew signal output
rlabel metal2 s 14830 49200 14886 50000 6 c_wb_o_dat[7]
port 59 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 c_wb_o_dat[8]
port 60 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 c_wb_o_dat[9]
port 61 nsew signal output
rlabel metal2 s 30930 49200 30986 50000 6 c_wb_sel[0]
port 62 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 c_wb_sel[1]
port 63 nsew signal output
rlabel metal3 s 39200 38768 40000 38888 6 c_wb_stb
port 64 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 c_wb_we
port 65 nsew signal output
rlabel metal3 s 39200 22448 40000 22568 6 cc_wb_4_burst
port 66 nsew signal input
rlabel metal2 s 10966 49200 11022 50000 6 cc_wb_8_burst
port 67 nsew signal input
rlabel metal2 s 38014 49200 38070 50000 6 cc_wb_adr[0]
port 68 nsew signal input
rlabel metal2 s 1950 49200 2006 50000 6 cc_wb_adr[10]
port 69 nsew signal input
rlabel metal3 s 39200 28568 40000 28688 6 cc_wb_adr[11]
port 70 nsew signal input
rlabel metal2 s 14186 49200 14242 50000 6 cc_wb_adr[12]
port 71 nsew signal input
rlabel metal3 s 39200 12248 40000 12368 6 cc_wb_adr[13]
port 72 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 cc_wb_adr[14]
port 73 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 cc_wb_adr[15]
port 74 nsew signal input
rlabel metal3 s 39200 17688 40000 17808 6 cc_wb_adr[16]
port 75 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 cc_wb_adr[17]
port 76 nsew signal input
rlabel metal3 s 39200 4088 40000 4208 6 cc_wb_adr[18]
port 77 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 cc_wb_adr[19]
port 78 nsew signal input
rlabel metal3 s 39200 11568 40000 11688 6 cc_wb_adr[1]
port 79 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 cc_wb_adr[20]
port 80 nsew signal input
rlabel metal3 s 39200 25168 40000 25288 6 cc_wb_adr[21]
port 81 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 cc_wb_adr[22]
port 82 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 cc_wb_adr[23]
port 83 nsew signal input
rlabel metal3 s 39200 10208 40000 10328 6 cc_wb_adr[2]
port 84 nsew signal input
rlabel metal3 s 39200 40808 40000 40928 6 cc_wb_adr[3]
port 85 nsew signal input
rlabel metal2 s 33506 49200 33562 50000 6 cc_wb_adr[4]
port 86 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 cc_wb_adr[5]
port 87 nsew signal input
rlabel metal3 s 39200 32648 40000 32768 6 cc_wb_adr[6]
port 88 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 cc_wb_adr[7]
port 89 nsew signal input
rlabel metal2 s 18694 49200 18750 50000 6 cc_wb_adr[8]
port 90 nsew signal input
rlabel metal3 s 39200 8 40000 128 6 cc_wb_adr[9]
port 91 nsew signal input
rlabel metal2 s 29642 49200 29698 50000 6 cc_wb_cyc
port 92 nsew signal input
rlabel metal3 s 39200 40128 40000 40248 6 cc_wb_o_dat[0]
port 93 nsew signal input
rlabel metal2 s 19338 49200 19394 50000 6 cc_wb_o_dat[10]
port 94 nsew signal input
rlabel metal2 s 5814 49200 5870 50000 6 cc_wb_o_dat[11]
port 95 nsew signal input
rlabel metal2 s 12898 49200 12954 50000 6 cc_wb_o_dat[12]
port 96 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 cc_wb_o_dat[13]
port 97 nsew signal input
rlabel metal2 s 23202 49200 23258 50000 6 cc_wb_o_dat[14]
port 98 nsew signal input
rlabel metal3 s 39200 17008 40000 17128 6 cc_wb_o_dat[15]
port 99 nsew signal input
rlabel metal3 s 39200 34008 40000 34128 6 cc_wb_o_dat[1]
port 100 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 cc_wb_o_dat[2]
port 101 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 cc_wb_o_dat[3]
port 102 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 cc_wb_o_dat[4]
port 103 nsew signal input
rlabel metal3 s 39200 46928 40000 47048 6 cc_wb_o_dat[5]
port 104 nsew signal input
rlabel metal3 s 0 688 800 808 6 cc_wb_o_dat[6]
port 105 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 cc_wb_o_dat[7]
port 106 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 cc_wb_o_dat[8]
port 107 nsew signal input
rlabel metal2 s 19982 49200 20038 50000 6 cc_wb_o_dat[9]
port 108 nsew signal input
rlabel metal2 s 16118 49200 16174 50000 6 cc_wb_sel[0]
port 109 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 cc_wb_sel[1]
port 110 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 cc_wb_stb
port 111 nsew signal input
rlabel metal2 s 39302 49200 39358 50000 6 cc_wb_we
port 112 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 cw_ack
port 113 nsew signal input
rlabel metal2 s 32862 49200 32918 50000 6 cw_clk
port 114 nsew signal input
rlabel metal2 s 21270 49200 21326 50000 6 cw_err
port 115 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 cw_io_i[0]
port 116 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 cw_io_i[10]
port 117 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 cw_io_i[11]
port 118 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 cw_io_i[12]
port 119 nsew signal input
rlabel metal2 s 18050 49200 18106 50000 6 cw_io_i[13]
port 120 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 cw_io_i[14]
port 121 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 cw_io_i[15]
port 122 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 cw_io_i[1]
port 123 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 cw_io_i[2]
port 124 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 cw_io_i[3]
port 125 nsew signal input
rlabel metal3 s 39200 29248 40000 29368 6 cw_io_i[4]
port 126 nsew signal input
rlabel metal2 s 38658 49200 38714 50000 6 cw_io_i[5]
port 127 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 cw_io_i[6]
port 128 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 cw_io_i[7]
port 129 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 cw_io_i[8]
port 130 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 cw_io_i[9]
port 131 nsew signal input
rlabel metal2 s 31574 49200 31630 50000 6 cw_rst
port 132 nsew signal output
rlabel metal3 s 39200 48288 40000 48408 6 cw_rst_z
port 133 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 i_clk
port 134 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 i_irq
port 135 nsew signal input
rlabel metal2 s 13542 49200 13598 50000 6 i_rst
port 136 nsew signal input
rlabel metal3 s 39200 9528 40000 9648 6 ic_split_clock
port 137 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 irq_s
port 138 nsew signal output
rlabel metal3 s 39200 30608 40000 30728 6 la_cw_ack
port 139 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_cw_io_i[0]
port 140 nsew signal input
rlabel metal3 s 39200 42168 40000 42288 6 la_cw_io_i[10]
port 141 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_cw_io_i[11]
port 142 nsew signal input
rlabel metal2 s 18 49200 74 50000 6 la_cw_io_i[12]
port 143 nsew signal input
rlabel metal2 s 9034 49200 9090 50000 6 la_cw_io_i[13]
port 144 nsew signal input
rlabel metal3 s 39200 10888 40000 11008 6 la_cw_io_i[14]
port 145 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 la_cw_io_i[15]
port 146 nsew signal input
rlabel metal3 s 39200 16328 40000 16448 6 la_cw_io_i[1]
port 147 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 la_cw_io_i[2]
port 148 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_cw_io_i[3]
port 149 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 la_cw_io_i[4]
port 150 nsew signal input
rlabel metal2 s 7102 49200 7158 50000 6 la_cw_io_i[5]
port 151 nsew signal input
rlabel metal3 s 39200 21768 40000 21888 6 la_cw_io_i[6]
port 152 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 la_cw_io_i[7]
port 153 nsew signal input
rlabel metal2 s 34794 49200 34850 50000 6 la_cw_io_i[8]
port 154 nsew signal input
rlabel metal3 s 39200 688 40000 808 6 la_cw_io_i[9]
port 155 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 la_cw_ovr
port 156 nsew signal input
rlabel metal3 s 39200 7488 40000 7608 6 m_cw_ack
port 157 nsew signal output
rlabel metal3 s 39200 44208 40000 44328 6 m_cw_err
port 158 nsew signal output
rlabel metal2 s 37370 49200 37426 50000 6 m_cw_io_i[0]
port 159 nsew signal output
rlabel metal2 s 22558 49200 22614 50000 6 m_cw_io_i[10]
port 160 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 m_cw_io_i[11]
port 161 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 m_cw_io_i[12]
port 162 nsew signal output
rlabel metal3 s 39200 23128 40000 23248 6 m_cw_io_i[13]
port 163 nsew signal output
rlabel metal3 s 39200 21088 40000 21208 6 m_cw_io_i[14]
port 164 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 m_cw_io_i[15]
port 165 nsew signal output
rlabel metal3 s 39200 18368 40000 18488 6 m_cw_io_i[1]
port 166 nsew signal output
rlabel metal3 s 39200 8168 40000 8288 6 m_cw_io_i[2]
port 167 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 m_cw_io_i[3]
port 168 nsew signal output
rlabel metal3 s 39200 47608 40000 47728 6 m_cw_io_i[4]
port 169 nsew signal output
rlabel metal3 s 39200 37408 40000 37528 6 m_cw_io_i[5]
port 170 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 m_cw_io_i[6]
port 171 nsew signal output
rlabel metal2 s 4526 49200 4582 50000 6 m_cw_io_i[7]
port 172 nsew signal output
rlabel metal3 s 39200 5448 40000 5568 6 m_cw_io_i[8]
port 173 nsew signal output
rlabel metal2 s 20626 49200 20682 50000 6 m_cw_io_i[9]
port 174 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 s_rst
port 175 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 u_wb_4_burst
port 176 nsew signal input
rlabel metal2 s 28354 49200 28410 50000 6 u_wb_8_burst
port 177 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 u_wb_ack
port 178 nsew signal output
rlabel metal3 s 39200 35368 40000 35488 6 u_wb_ack_cc
port 179 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 u_wb_ack_clk
port 180 nsew signal output
rlabel metal3 s 39200 44888 40000 45008 6 u_wb_ack_mxed
port 181 nsew signal output
rlabel metal3 s 39200 14288 40000 14408 6 u_wb_adr[0]
port 182 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 u_wb_adr[10]
port 183 nsew signal input
rlabel metal3 s 39200 46248 40000 46368 6 u_wb_adr[11]
port 184 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 u_wb_adr[12]
port 185 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 u_wb_adr[13]
port 186 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 u_wb_adr[14]
port 187 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 u_wb_adr[15]
port 188 nsew signal input
rlabel metal3 s 39200 8848 40000 8968 6 u_wb_adr[16]
port 189 nsew signal input
rlabel metal2 s 23846 49200 23902 50000 6 u_wb_adr[17]
port 190 nsew signal input
rlabel metal3 s 39200 33328 40000 33448 6 u_wb_adr[18]
port 191 nsew signal input
rlabel metal2 s 2594 49200 2650 50000 6 u_wb_adr[19]
port 192 nsew signal input
rlabel metal2 s 5170 49200 5226 50000 6 u_wb_adr[1]
port 193 nsew signal input
rlabel metal2 s 3238 49200 3294 50000 6 u_wb_adr[20]
port 194 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 u_wb_adr[21]
port 195 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 u_wb_adr[22]
port 196 nsew signal input
rlabel metal3 s 39200 20408 40000 20528 6 u_wb_adr[23]
port 197 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 u_wb_adr[2]
port 198 nsew signal input
rlabel metal2 s 36082 49200 36138 50000 6 u_wb_adr[3]
port 199 nsew signal input
rlabel metal3 s 39200 43528 40000 43648 6 u_wb_adr[4]
port 200 nsew signal input
rlabel metal2 s 11610 49200 11666 50000 6 u_wb_adr[5]
port 201 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 u_wb_adr[6]
port 202 nsew signal input
rlabel metal3 s 39200 24488 40000 24608 6 u_wb_adr[7]
port 203 nsew signal input
rlabel metal3 s 39200 42848 40000 42968 6 u_wb_adr[8]
port 204 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 u_wb_adr[9]
port 205 nsew signal input
rlabel metal3 s 39200 31968 40000 32088 6 u_wb_cyc
port 206 nsew signal input
rlabel metal3 s 39200 13608 40000 13728 6 u_wb_err
port 207 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 u_wb_err_cc
port 208 nsew signal input
rlabel metal3 s 39200 48968 40000 49088 6 u_wb_i_dat[0]
port 209 nsew signal output
rlabel metal2 s 16762 49200 16818 50000 6 u_wb_i_dat[10]
port 210 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 u_wb_i_dat[11]
port 211 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 u_wb_i_dat[12]
port 212 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 u_wb_i_dat[13]
port 213 nsew signal output
rlabel metal3 s 39200 12928 40000 13048 6 u_wb_i_dat[14]
port 214 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 u_wb_i_dat[15]
port 215 nsew signal output
rlabel metal3 s 39200 2048 40000 2168 6 u_wb_i_dat[1]
port 216 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 u_wb_i_dat[2]
port 217 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 u_wb_i_dat[3]
port 218 nsew signal output
rlabel metal3 s 39200 19728 40000 19848 6 u_wb_i_dat[4]
port 219 nsew signal output
rlabel metal2 s 36726 49200 36782 50000 6 u_wb_i_dat[5]
port 220 nsew signal output
rlabel metal3 s 39200 39448 40000 39568 6 u_wb_i_dat[6]
port 221 nsew signal output
rlabel metal3 s 39200 2728 40000 2848 6 u_wb_i_dat[7]
port 222 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 u_wb_i_dat[8]
port 223 nsew signal output
rlabel metal3 s 39200 25848 40000 25968 6 u_wb_i_dat[9]
port 224 nsew signal output
rlabel metal2 s 662 0 718 800 6 u_wb_i_dat_cc[0]
port 225 nsew signal input
rlabel metal3 s 39200 41488 40000 41608 6 u_wb_i_dat_cc[10]
port 226 nsew signal input
rlabel metal2 s 34150 49200 34206 50000 6 u_wb_i_dat_cc[11]
port 227 nsew signal input
rlabel metal3 s 39200 6808 40000 6928 6 u_wb_i_dat_cc[12]
port 228 nsew signal input
rlabel metal2 s 32218 49200 32274 50000 6 u_wb_i_dat_cc[13]
port 229 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 u_wb_i_dat_cc[14]
port 230 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 u_wb_i_dat_cc[15]
port 231 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 u_wb_i_dat_cc[1]
port 232 nsew signal input
rlabel metal2 s 18 0 74 800 6 u_wb_i_dat_cc[2]
port 233 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 u_wb_i_dat_cc[3]
port 234 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 u_wb_i_dat_cc[4]
port 235 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 u_wb_i_dat_cc[5]
port 236 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 u_wb_i_dat_cc[6]
port 237 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 u_wb_i_dat_cc[7]
port 238 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 u_wb_i_dat_cc[8]
port 239 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 u_wb_i_dat_cc[9]
port 240 nsew signal input
rlabel metal2 s 21914 49200 21970 50000 6 u_wb_o_dat[0]
port 241 nsew signal input
rlabel metal2 s 12254 49200 12310 50000 6 u_wb_o_dat[10]
port 242 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 u_wb_o_dat[11]
port 243 nsew signal input
rlabel metal2 s 28998 49200 29054 50000 6 u_wb_o_dat[12]
port 244 nsew signal input
rlabel metal3 s 39200 14968 40000 15088 6 u_wb_o_dat[13]
port 245 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 u_wb_o_dat[14]
port 246 nsew signal input
rlabel metal3 s 39200 38088 40000 38208 6 u_wb_o_dat[15]
port 247 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 u_wb_o_dat[1]
port 248 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 u_wb_o_dat[2]
port 249 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 u_wb_o_dat[3]
port 250 nsew signal input
rlabel metal3 s 39200 36728 40000 36848 6 u_wb_o_dat[4]
port 251 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 u_wb_o_dat[5]
port 252 nsew signal input
rlabel metal2 s 25778 49200 25834 50000 6 u_wb_o_dat[6]
port 253 nsew signal input
rlabel metal2 s 24490 49200 24546 50000 6 u_wb_o_dat[7]
port 254 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 u_wb_o_dat[8]
port 255 nsew signal input
rlabel metal2 s 1306 49200 1362 50000 6 u_wb_o_dat[9]
port 256 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 u_wb_sel[0]
port 257 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 u_wb_sel[1]
port 258 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 u_wb_stb
port 259 nsew signal input
rlabel metal3 s 39200 26528 40000 26648 6 u_wb_we
port 260 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 261 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 261 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 262 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1770760
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/top_cw_logic/runs/22_09_13_13_56/results/signoff/top_cw_logic.magic.gds
string GDS_START 183926
<< end >>

