magic
tech gf180mcuD
timestamp 1700048757
<< metal5 >>
rect 0 1400 400 1600
rect 1000 1400 1400 1600
rect 8800 1400 10220 1600
rect 0 400 200 1400
rect 580 780 820 1020
rect 600 600 660 620
rect 580 580 720 600
rect 580 560 780 580
rect 580 540 820 560
rect 560 480 820 540
rect 540 420 800 480
rect 0 360 400 400
rect 520 360 780 420
rect 1200 400 1400 1400
rect 9080 1320 9280 1400
rect 9060 1300 9280 1320
rect 9720 1300 9920 1400
rect 9060 1220 9260 1300
rect 9040 1200 9260 1220
rect 9700 1200 9900 1300
rect 9040 1120 9240 1200
rect 9020 1100 9240 1120
rect 9680 1100 9880 1200
rect 12800 1100 13200 1200
rect 5700 1020 6000 1100
rect 6620 1040 6800 1100
rect 6560 1020 6800 1040
rect 5700 1000 6020 1020
rect 1000 360 1400 400
rect 0 320 380 360
rect 0 260 360 320
rect 500 300 760 360
rect 980 320 1400 360
rect 480 260 740 300
rect 960 260 1400 320
rect 0 200 340 260
rect 480 240 720 260
rect 460 200 720 240
rect 940 200 1400 260
rect 1700 820 2200 900
rect 2500 820 2900 900
rect 3300 820 3700 900
rect 1700 800 2220 820
rect 2500 800 2920 820
rect 3280 800 3700 820
rect 3800 820 4200 900
rect 3800 800 4220 820
rect 1700 500 1900 800
rect 2180 780 2300 800
rect 2200 520 2300 780
rect 2180 500 2300 520
rect 2500 500 2600 800
rect 2880 780 3000 800
rect 2900 520 3000 780
rect 2880 500 3000 520
rect 3200 780 3320 800
rect 3200 520 3300 780
rect 3200 500 3320 520
rect 3800 500 3900 800
rect 4180 780 4300 800
rect 4200 520 4300 780
rect 4180 500 4300 520
rect 4400 520 4500 860
rect 4800 520 4900 860
rect 6000 820 6100 1000
rect 6560 980 6640 1020
rect 6500 960 6640 980
rect 6500 920 6580 960
rect 6440 900 6580 920
rect 6440 860 6520 900
rect 6400 840 6520 860
rect 6400 820 6460 840
rect 5980 800 6100 820
rect 6380 800 6460 820
rect 5700 720 6000 800
rect 6340 780 6460 800
rect 6340 760 6440 780
rect 6700 760 6800 1020
rect 7100 900 7200 1040
rect 7500 1020 7800 1100
rect 7480 1000 7820 1020
rect 9020 1000 9220 1100
rect 9660 1000 9860 1100
rect 10600 1020 10900 1100
rect 10580 1000 10900 1020
rect 11000 1000 11400 1100
rect 6960 800 7340 900
rect 7400 800 7500 1000
rect 7800 800 7900 1000
rect 9000 900 9200 1000
rect 9640 900 9840 1000
rect 10500 980 10640 1000
rect 11260 980 11400 1000
rect 10500 960 10620 980
rect 11280 960 11400 980
rect 10500 940 10600 960
rect 10500 920 10620 940
rect 11300 920 11400 960
rect 10500 900 10640 920
rect 11280 900 11400 920
rect 11500 1000 11900 1100
rect 12000 1000 12400 1100
rect 11500 980 11620 1000
rect 12000 980 12120 1000
rect 11500 920 11600 980
rect 12000 920 12100 980
rect 11500 900 11620 920
rect 12000 900 12120 920
rect 13100 900 13200 1100
rect 8980 800 9180 900
rect 9620 800 9820 900
rect 10600 840 10800 900
rect 11240 880 11360 900
rect 11220 860 11340 880
rect 11200 840 11320 860
rect 10600 820 10820 840
rect 11180 820 11300 840
rect 10600 800 10840 820
rect 11160 800 11280 820
rect 11500 800 11900 900
rect 12000 800 12400 900
rect 12800 800 13200 900
rect 13300 1100 13800 1200
rect 13900 1100 14300 1200
rect 14400 1100 14800 1200
rect 6340 720 6800 760
rect 5700 700 6020 720
rect 6360 700 6800 720
rect 5980 680 6100 700
rect 4400 500 4520 520
rect 4780 500 4900 520
rect 6000 500 6100 680
rect 6380 660 6800 700
rect 7100 660 7200 800
rect 7460 780 7840 800
rect 7480 760 7820 780
rect 7500 740 7800 760
rect 7480 720 7820 740
rect 7460 700 7840 720
rect 8960 700 9160 800
rect 9600 700 9800 800
rect 10780 780 10900 800
rect 11140 780 11260 800
rect 11500 780 11620 800
rect 1700 480 2220 500
rect 2500 480 2920 500
rect 3280 480 3700 500
rect 1700 400 2200 480
rect 2500 400 2900 480
rect 3300 400 3700 480
rect 3800 480 4220 500
rect 4480 480 4800 500
rect 3800 400 4200 480
rect 4500 400 4800 480
rect 5700 480 6020 500
rect 5700 400 6000 480
rect 6200 400 6300 500
rect 6700 400 6800 660
rect 6980 500 7320 600
rect 7400 500 7500 700
rect 7800 500 7900 700
rect 8940 600 9140 700
rect 9580 640 9800 700
rect 9580 600 9880 640
rect 10800 620 10900 780
rect 11120 760 11240 780
rect 11100 740 11220 760
rect 11080 720 11200 740
rect 11060 700 11180 720
rect 11020 680 11160 700
rect 10780 600 10900 620
rect 11000 660 11140 680
rect 11000 640 11120 660
rect 11000 620 11100 640
rect 11500 620 11600 780
rect 11000 600 11120 620
rect 11500 600 11620 620
rect 8920 500 9120 600
rect 9560 560 9880 600
rect 10500 580 10840 600
rect 10500 560 10820 580
rect 9560 500 9860 560
rect 10500 500 10800 560
rect 11000 500 11400 600
rect 11500 500 11900 600
rect 12000 500 12100 800
rect 12800 600 12900 800
rect 13300 600 13400 1100
rect 13700 600 13800 1100
rect 14200 900 14300 1100
rect 14700 900 14800 1100
rect 12800 500 13200 600
rect 13300 500 13800 600
rect 13900 800 14300 900
rect 14400 800 14800 900
rect 13900 600 14000 800
rect 14700 600 14800 800
rect 13900 500 14300 600
rect 14400 500 14800 600
rect 7480 480 7820 500
rect 7500 400 7800 480
rect 480 180 700 200
rect 560 160 700 180
rect 620 140 700 160
rect 1700 0 1900 400
rect 2500 0 2600 400
rect 3800 0 3900 400
<< end >>
