VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO icache
  CLASS BLOCK ;
  FOREIGN icache ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 1770.000 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.360 4.000 59.920 ;
    END
  END i_clk
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.280 4.000 77.840 ;
    END
  END i_rst
  PIN mem_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.200 4.000 95.760 ;
    END
  END mem_ack
  PIN mem_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 256.480 4.000 257.040 ;
    END
  END mem_addr[0]
  PIN mem_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1009.120 4.000 1009.680 ;
    END
  END mem_addr[10]
  PIN mem_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1080.800 4.000 1081.360 ;
    END
  END mem_addr[11]
  PIN mem_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1152.480 4.000 1153.040 ;
    END
  END mem_addr[12]
  PIN mem_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1224.160 4.000 1224.720 ;
    END
  END mem_addr[13]
  PIN mem_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1295.840 4.000 1296.400 ;
    END
  END mem_addr[14]
  PIN mem_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1367.520 4.000 1368.080 ;
    END
  END mem_addr[15]
  PIN mem_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 346.080 4.000 346.640 ;
    END
  END mem_addr[1]
  PIN mem_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 435.680 4.000 436.240 ;
    END
  END mem_addr[2]
  PIN mem_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 507.360 4.000 507.920 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 579.040 4.000 579.600 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 650.720 4.000 651.280 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 722.400 4.000 722.960 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 794.080 4.000 794.640 ;
    END
  END mem_addr[7]
  PIN mem_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 865.760 4.000 866.320 ;
    END
  END mem_addr[8]
  PIN mem_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 937.440 4.000 938.000 ;
    END
  END mem_addr[9]
  PIN mem_cache_flush
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 113.120 4.000 113.680 ;
    END
  END mem_cache_flush
  PIN mem_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 274.400 4.000 274.960 ;
    END
  END mem_data[0]
  PIN mem_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1027.040 4.000 1027.600 ;
    END
  END mem_data[10]
  PIN mem_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1098.720 4.000 1099.280 ;
    END
  END mem_data[11]
  PIN mem_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1170.400 4.000 1170.960 ;
    END
  END mem_data[12]
  PIN mem_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1242.080 4.000 1242.640 ;
    END
  END mem_data[13]
  PIN mem_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1313.760 4.000 1314.320 ;
    END
  END mem_data[14]
  PIN mem_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1385.440 4.000 1386.000 ;
    END
  END mem_data[15]
  PIN mem_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1439.200 4.000 1439.760 ;
    END
  END mem_data[16]
  PIN mem_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1457.120 4.000 1457.680 ;
    END
  END mem_data[17]
  PIN mem_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1475.040 4.000 1475.600 ;
    END
  END mem_data[18]
  PIN mem_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1492.960 4.000 1493.520 ;
    END
  END mem_data[19]
  PIN mem_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 364.000 4.000 364.560 ;
    END
  END mem_data[1]
  PIN mem_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1510.880 4.000 1511.440 ;
    END
  END mem_data[20]
  PIN mem_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1528.800 4.000 1529.360 ;
    END
  END mem_data[21]
  PIN mem_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1546.720 4.000 1547.280 ;
    END
  END mem_data[22]
  PIN mem_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1564.640 4.000 1565.200 ;
    END
  END mem_data[23]
  PIN mem_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1582.560 4.000 1583.120 ;
    END
  END mem_data[24]
  PIN mem_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1600.480 4.000 1601.040 ;
    END
  END mem_data[25]
  PIN mem_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1618.400 4.000 1618.960 ;
    END
  END mem_data[26]
  PIN mem_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1636.320 4.000 1636.880 ;
    END
  END mem_data[27]
  PIN mem_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1654.240 4.000 1654.800 ;
    END
  END mem_data[28]
  PIN mem_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1672.160 4.000 1672.720 ;
    END
  END mem_data[29]
  PIN mem_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 453.600 4.000 454.160 ;
    END
  END mem_data[2]
  PIN mem_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1690.080 4.000 1690.640 ;
    END
  END mem_data[30]
  PIN mem_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1708.000 4.000 1708.560 ;
    END
  END mem_data[31]
  PIN mem_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 525.280 4.000 525.840 ;
    END
  END mem_data[3]
  PIN mem_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 596.960 4.000 597.520 ;
    END
  END mem_data[4]
  PIN mem_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 668.640 4.000 669.200 ;
    END
  END mem_data[5]
  PIN mem_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 740.320 4.000 740.880 ;
    END
  END mem_data[6]
  PIN mem_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 812.000 4.000 812.560 ;
    END
  END mem_data[7]
  PIN mem_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 883.680 4.000 884.240 ;
    END
  END mem_data[8]
  PIN mem_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 955.360 4.000 955.920 ;
    END
  END mem_data[9]
  PIN mem_ppl_submit
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END mem_ppl_submit
  PIN mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 148.960 4.000 149.520 ;
    END
  END mem_req
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1752.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1752.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1752.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1752.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1752.540 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1752.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1752.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1752.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1752.540 ;
    END
  END vssd1
  PIN wb_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.880 4.000 167.440 ;
    END
  END wb_ack
  PIN wb_adr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 292.320 4.000 292.880 ;
    END
  END wb_adr[0]
  PIN wb_adr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1044.960 4.000 1045.520 ;
    END
  END wb_adr[10]
  PIN wb_adr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1116.640 4.000 1117.200 ;
    END
  END wb_adr[11]
  PIN wb_adr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1188.320 4.000 1188.880 ;
    END
  END wb_adr[12]
  PIN wb_adr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1260.000 4.000 1260.560 ;
    END
  END wb_adr[13]
  PIN wb_adr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1331.680 4.000 1332.240 ;
    END
  END wb_adr[14]
  PIN wb_adr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1403.360 4.000 1403.920 ;
    END
  END wb_adr[15]
  PIN wb_adr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 381.920 4.000 382.480 ;
    END
  END wb_adr[1]
  PIN wb_adr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 471.520 4.000 472.080 ;
    END
  END wb_adr[2]
  PIN wb_adr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 543.200 4.000 543.760 ;
    END
  END wb_adr[3]
  PIN wb_adr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 614.880 4.000 615.440 ;
    END
  END wb_adr[4]
  PIN wb_adr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 686.560 4.000 687.120 ;
    END
  END wb_adr[5]
  PIN wb_adr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 758.240 4.000 758.800 ;
    END
  END wb_adr[6]
  PIN wb_adr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 829.920 4.000 830.480 ;
    END
  END wb_adr[7]
  PIN wb_adr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 901.600 4.000 902.160 ;
    END
  END wb_adr[8]
  PIN wb_adr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 973.280 4.000 973.840 ;
    END
  END wb_adr[9]
  PIN wb_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END wb_cyc
  PIN wb_err
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 202.720 4.000 203.280 ;
    END
  END wb_err
  PIN wb_i_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.240 4.000 310.800 ;
    END
  END wb_i_dat[0]
  PIN wb_i_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1062.880 4.000 1063.440 ;
    END
  END wb_i_dat[10]
  PIN wb_i_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1134.560 4.000 1135.120 ;
    END
  END wb_i_dat[11]
  PIN wb_i_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1206.240 4.000 1206.800 ;
    END
  END wb_i_dat[12]
  PIN wb_i_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1277.920 4.000 1278.480 ;
    END
  END wb_i_dat[13]
  PIN wb_i_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1349.600 4.000 1350.160 ;
    END
  END wb_i_dat[14]
  PIN wb_i_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1421.280 4.000 1421.840 ;
    END
  END wb_i_dat[15]
  PIN wb_i_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 399.840 4.000 400.400 ;
    END
  END wb_i_dat[1]
  PIN wb_i_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 489.440 4.000 490.000 ;
    END
  END wb_i_dat[2]
  PIN wb_i_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 561.120 4.000 561.680 ;
    END
  END wb_i_dat[3]
  PIN wb_i_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 632.800 4.000 633.360 ;
    END
  END wb_i_dat[4]
  PIN wb_i_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 704.480 4.000 705.040 ;
    END
  END wb_i_dat[5]
  PIN wb_i_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 776.160 4.000 776.720 ;
    END
  END wb_i_dat[6]
  PIN wb_i_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 847.840 4.000 848.400 ;
    END
  END wb_i_dat[7]
  PIN wb_i_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 919.520 4.000 920.080 ;
    END
  END wb_i_dat[8]
  PIN wb_i_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 991.200 4.000 991.760 ;
    END
  END wb_i_dat[9]
  PIN wb_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 328.160 4.000 328.720 ;
    END
  END wb_sel[0]
  PIN wb_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 417.760 4.000 418.320 ;
    END
  END wb_sel[1]
  PIN wb_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 220.640 4.000 221.200 ;
    END
  END wb_stb
  PIN wb_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 4.000 239.120 ;
    END
  END wb_we
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 693.280 1752.540 ;
      LAYER Metal2 ;
        RECT 1.820 5.690 694.260 1752.430 ;
      LAYER Metal3 ;
        RECT 1.770 1708.860 694.310 1752.380 ;
        RECT 4.300 1707.700 694.310 1708.860 ;
        RECT 1.770 1690.940 694.310 1707.700 ;
        RECT 4.300 1689.780 694.310 1690.940 ;
        RECT 1.770 1673.020 694.310 1689.780 ;
        RECT 4.300 1671.860 694.310 1673.020 ;
        RECT 1.770 1655.100 694.310 1671.860 ;
        RECT 4.300 1653.940 694.310 1655.100 ;
        RECT 1.770 1637.180 694.310 1653.940 ;
        RECT 4.300 1636.020 694.310 1637.180 ;
        RECT 1.770 1619.260 694.310 1636.020 ;
        RECT 4.300 1618.100 694.310 1619.260 ;
        RECT 1.770 1601.340 694.310 1618.100 ;
        RECT 4.300 1600.180 694.310 1601.340 ;
        RECT 1.770 1583.420 694.310 1600.180 ;
        RECT 4.300 1582.260 694.310 1583.420 ;
        RECT 1.770 1565.500 694.310 1582.260 ;
        RECT 4.300 1564.340 694.310 1565.500 ;
        RECT 1.770 1547.580 694.310 1564.340 ;
        RECT 4.300 1546.420 694.310 1547.580 ;
        RECT 1.770 1529.660 694.310 1546.420 ;
        RECT 4.300 1528.500 694.310 1529.660 ;
        RECT 1.770 1511.740 694.310 1528.500 ;
        RECT 4.300 1510.580 694.310 1511.740 ;
        RECT 1.770 1493.820 694.310 1510.580 ;
        RECT 4.300 1492.660 694.310 1493.820 ;
        RECT 1.770 1475.900 694.310 1492.660 ;
        RECT 4.300 1474.740 694.310 1475.900 ;
        RECT 1.770 1457.980 694.310 1474.740 ;
        RECT 4.300 1456.820 694.310 1457.980 ;
        RECT 1.770 1440.060 694.310 1456.820 ;
        RECT 4.300 1438.900 694.310 1440.060 ;
        RECT 1.770 1422.140 694.310 1438.900 ;
        RECT 4.300 1420.980 694.310 1422.140 ;
        RECT 1.770 1404.220 694.310 1420.980 ;
        RECT 4.300 1403.060 694.310 1404.220 ;
        RECT 1.770 1386.300 694.310 1403.060 ;
        RECT 4.300 1385.140 694.310 1386.300 ;
        RECT 1.770 1368.380 694.310 1385.140 ;
        RECT 4.300 1367.220 694.310 1368.380 ;
        RECT 1.770 1350.460 694.310 1367.220 ;
        RECT 4.300 1349.300 694.310 1350.460 ;
        RECT 1.770 1332.540 694.310 1349.300 ;
        RECT 4.300 1331.380 694.310 1332.540 ;
        RECT 1.770 1314.620 694.310 1331.380 ;
        RECT 4.300 1313.460 694.310 1314.620 ;
        RECT 1.770 1296.700 694.310 1313.460 ;
        RECT 4.300 1295.540 694.310 1296.700 ;
        RECT 1.770 1278.780 694.310 1295.540 ;
        RECT 4.300 1277.620 694.310 1278.780 ;
        RECT 1.770 1260.860 694.310 1277.620 ;
        RECT 4.300 1259.700 694.310 1260.860 ;
        RECT 1.770 1242.940 694.310 1259.700 ;
        RECT 4.300 1241.780 694.310 1242.940 ;
        RECT 1.770 1225.020 694.310 1241.780 ;
        RECT 4.300 1223.860 694.310 1225.020 ;
        RECT 1.770 1207.100 694.310 1223.860 ;
        RECT 4.300 1205.940 694.310 1207.100 ;
        RECT 1.770 1189.180 694.310 1205.940 ;
        RECT 4.300 1188.020 694.310 1189.180 ;
        RECT 1.770 1171.260 694.310 1188.020 ;
        RECT 4.300 1170.100 694.310 1171.260 ;
        RECT 1.770 1153.340 694.310 1170.100 ;
        RECT 4.300 1152.180 694.310 1153.340 ;
        RECT 1.770 1135.420 694.310 1152.180 ;
        RECT 4.300 1134.260 694.310 1135.420 ;
        RECT 1.770 1117.500 694.310 1134.260 ;
        RECT 4.300 1116.340 694.310 1117.500 ;
        RECT 1.770 1099.580 694.310 1116.340 ;
        RECT 4.300 1098.420 694.310 1099.580 ;
        RECT 1.770 1081.660 694.310 1098.420 ;
        RECT 4.300 1080.500 694.310 1081.660 ;
        RECT 1.770 1063.740 694.310 1080.500 ;
        RECT 4.300 1062.580 694.310 1063.740 ;
        RECT 1.770 1045.820 694.310 1062.580 ;
        RECT 4.300 1044.660 694.310 1045.820 ;
        RECT 1.770 1027.900 694.310 1044.660 ;
        RECT 4.300 1026.740 694.310 1027.900 ;
        RECT 1.770 1009.980 694.310 1026.740 ;
        RECT 4.300 1008.820 694.310 1009.980 ;
        RECT 1.770 992.060 694.310 1008.820 ;
        RECT 4.300 990.900 694.310 992.060 ;
        RECT 1.770 974.140 694.310 990.900 ;
        RECT 4.300 972.980 694.310 974.140 ;
        RECT 1.770 956.220 694.310 972.980 ;
        RECT 4.300 955.060 694.310 956.220 ;
        RECT 1.770 938.300 694.310 955.060 ;
        RECT 4.300 937.140 694.310 938.300 ;
        RECT 1.770 920.380 694.310 937.140 ;
        RECT 4.300 919.220 694.310 920.380 ;
        RECT 1.770 902.460 694.310 919.220 ;
        RECT 4.300 901.300 694.310 902.460 ;
        RECT 1.770 884.540 694.310 901.300 ;
        RECT 4.300 883.380 694.310 884.540 ;
        RECT 1.770 866.620 694.310 883.380 ;
        RECT 4.300 865.460 694.310 866.620 ;
        RECT 1.770 848.700 694.310 865.460 ;
        RECT 4.300 847.540 694.310 848.700 ;
        RECT 1.770 830.780 694.310 847.540 ;
        RECT 4.300 829.620 694.310 830.780 ;
        RECT 1.770 812.860 694.310 829.620 ;
        RECT 4.300 811.700 694.310 812.860 ;
        RECT 1.770 794.940 694.310 811.700 ;
        RECT 4.300 793.780 694.310 794.940 ;
        RECT 1.770 777.020 694.310 793.780 ;
        RECT 4.300 775.860 694.310 777.020 ;
        RECT 1.770 759.100 694.310 775.860 ;
        RECT 4.300 757.940 694.310 759.100 ;
        RECT 1.770 741.180 694.310 757.940 ;
        RECT 4.300 740.020 694.310 741.180 ;
        RECT 1.770 723.260 694.310 740.020 ;
        RECT 4.300 722.100 694.310 723.260 ;
        RECT 1.770 705.340 694.310 722.100 ;
        RECT 4.300 704.180 694.310 705.340 ;
        RECT 1.770 687.420 694.310 704.180 ;
        RECT 4.300 686.260 694.310 687.420 ;
        RECT 1.770 669.500 694.310 686.260 ;
        RECT 4.300 668.340 694.310 669.500 ;
        RECT 1.770 651.580 694.310 668.340 ;
        RECT 4.300 650.420 694.310 651.580 ;
        RECT 1.770 633.660 694.310 650.420 ;
        RECT 4.300 632.500 694.310 633.660 ;
        RECT 1.770 615.740 694.310 632.500 ;
        RECT 4.300 614.580 694.310 615.740 ;
        RECT 1.770 597.820 694.310 614.580 ;
        RECT 4.300 596.660 694.310 597.820 ;
        RECT 1.770 579.900 694.310 596.660 ;
        RECT 4.300 578.740 694.310 579.900 ;
        RECT 1.770 561.980 694.310 578.740 ;
        RECT 4.300 560.820 694.310 561.980 ;
        RECT 1.770 544.060 694.310 560.820 ;
        RECT 4.300 542.900 694.310 544.060 ;
        RECT 1.770 526.140 694.310 542.900 ;
        RECT 4.300 524.980 694.310 526.140 ;
        RECT 1.770 508.220 694.310 524.980 ;
        RECT 4.300 507.060 694.310 508.220 ;
        RECT 1.770 490.300 694.310 507.060 ;
        RECT 4.300 489.140 694.310 490.300 ;
        RECT 1.770 472.380 694.310 489.140 ;
        RECT 4.300 471.220 694.310 472.380 ;
        RECT 1.770 454.460 694.310 471.220 ;
        RECT 4.300 453.300 694.310 454.460 ;
        RECT 1.770 436.540 694.310 453.300 ;
        RECT 4.300 435.380 694.310 436.540 ;
        RECT 1.770 418.620 694.310 435.380 ;
        RECT 4.300 417.460 694.310 418.620 ;
        RECT 1.770 400.700 694.310 417.460 ;
        RECT 4.300 399.540 694.310 400.700 ;
        RECT 1.770 382.780 694.310 399.540 ;
        RECT 4.300 381.620 694.310 382.780 ;
        RECT 1.770 364.860 694.310 381.620 ;
        RECT 4.300 363.700 694.310 364.860 ;
        RECT 1.770 346.940 694.310 363.700 ;
        RECT 4.300 345.780 694.310 346.940 ;
        RECT 1.770 329.020 694.310 345.780 ;
        RECT 4.300 327.860 694.310 329.020 ;
        RECT 1.770 311.100 694.310 327.860 ;
        RECT 4.300 309.940 694.310 311.100 ;
        RECT 1.770 293.180 694.310 309.940 ;
        RECT 4.300 292.020 694.310 293.180 ;
        RECT 1.770 275.260 694.310 292.020 ;
        RECT 4.300 274.100 694.310 275.260 ;
        RECT 1.770 257.340 694.310 274.100 ;
        RECT 4.300 256.180 694.310 257.340 ;
        RECT 1.770 239.420 694.310 256.180 ;
        RECT 4.300 238.260 694.310 239.420 ;
        RECT 1.770 221.500 694.310 238.260 ;
        RECT 4.300 220.340 694.310 221.500 ;
        RECT 1.770 203.580 694.310 220.340 ;
        RECT 4.300 202.420 694.310 203.580 ;
        RECT 1.770 185.660 694.310 202.420 ;
        RECT 4.300 184.500 694.310 185.660 ;
        RECT 1.770 167.740 694.310 184.500 ;
        RECT 4.300 166.580 694.310 167.740 ;
        RECT 1.770 149.820 694.310 166.580 ;
        RECT 4.300 148.660 694.310 149.820 ;
        RECT 1.770 131.900 694.310 148.660 ;
        RECT 4.300 130.740 694.310 131.900 ;
        RECT 1.770 113.980 694.310 130.740 ;
        RECT 4.300 112.820 694.310 113.980 ;
        RECT 1.770 96.060 694.310 112.820 ;
        RECT 4.300 94.900 694.310 96.060 ;
        RECT 1.770 78.140 694.310 94.900 ;
        RECT 4.300 76.980 694.310 78.140 ;
        RECT 1.770 60.220 694.310 76.980 ;
        RECT 4.300 59.060 694.310 60.220 ;
        RECT 1.770 5.740 694.310 59.060 ;
      LAYER Metal4 ;
        RECT 7.420 15.080 21.940 1749.910 ;
        RECT 24.140 15.080 98.740 1749.910 ;
        RECT 100.940 15.080 175.540 1749.910 ;
        RECT 177.740 15.080 252.340 1749.910 ;
        RECT 254.540 15.080 329.140 1749.910 ;
        RECT 331.340 15.080 405.940 1749.910 ;
        RECT 408.140 15.080 482.740 1749.910 ;
        RECT 484.940 15.080 559.540 1749.910 ;
        RECT 561.740 15.080 636.340 1749.910 ;
        RECT 638.540 15.080 691.460 1749.910 ;
        RECT 7.420 5.690 691.460 15.080 ;
  END
END icache
END LIBRARY

