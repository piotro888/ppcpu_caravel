// This is the unpowered netlist.
module core0 (i_clk,
    i_disable,
    i_irq,
    i_mc_core_int,
    i_mem_ack,
    i_mem_exception,
    i_req_data_valid,
    i_rst,
    o_c_data_page,
    o_c_instr_long,
    o_c_instr_page,
    o_icache_flush,
    o_mem_long,
    o_mem_req,
    o_mem_we,
    o_req_active,
    o_req_ppl_submit,
    sr_bus_we,
    dbg_pc,
    dbg_r0,
    i_core_int_sreg,
    i_mem_data,
    i_req_data,
    o_instr_long_addr,
    o_mem_addr,
    o_mem_addr_high,
    o_mem_data,
    o_mem_sel,
    o_req_addr,
    sr_bus_addr,
    sr_bus_data_o);
 input i_clk;
 input i_disable;
 input i_irq;
 input i_mc_core_int;
 input i_mem_ack;
 input i_mem_exception;
 input i_req_data_valid;
 input i_rst;
 output o_c_data_page;
 output o_c_instr_long;
 output o_c_instr_page;
 output o_icache_flush;
 output o_mem_long;
 output o_mem_req;
 output o_mem_we;
 output o_req_active;
 output o_req_ppl_submit;
 output sr_bus_we;
 output [15:0] dbg_pc;
 output [15:0] dbg_r0;
 input [15:0] i_core_int_sreg;
 input [15:0] i_mem_data;
 input [31:0] i_req_data;
 output [7:0] o_instr_long_addr;
 output [15:0] o_mem_addr;
 output [7:0] o_mem_addr_high;
 output [15:0] o_mem_data;
 output [1:0] o_mem_sel;
 output [15:0] o_req_addr;
 output [15:0] sr_bus_addr;
 output [15:0] sr_bus_data_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire \core_0.de_jmp_pred ;
 wire \core_0.dec_alu_carry_en ;
 wire \core_0.dec_alu_flags_ie ;
 wire \core_0.dec_jump_cond_code[0] ;
 wire \core_0.dec_jump_cond_code[1] ;
 wire \core_0.dec_jump_cond_code[2] ;
 wire \core_0.dec_jump_cond_code[3] ;
 wire \core_0.dec_jump_cond_code[4] ;
 wire \core_0.dec_l_reg_sel[0] ;
 wire \core_0.dec_l_reg_sel[1] ;
 wire \core_0.dec_l_reg_sel[2] ;
 wire \core_0.dec_mem_access ;
 wire \core_0.dec_mem_long ;
 wire \core_0.dec_mem_we ;
 wire \core_0.dec_mem_width ;
 wire \core_0.dec_pc_inc ;
 wire \core_0.dec_r_bus_imm ;
 wire \core_0.dec_r_reg_sel[0] ;
 wire \core_0.dec_r_reg_sel[1] ;
 wire \core_0.dec_r_reg_sel[2] ;
 wire \core_0.dec_rf_ie[0] ;
 wire \core_0.dec_rf_ie[1] ;
 wire \core_0.dec_rf_ie[2] ;
 wire \core_0.dec_rf_ie[3] ;
 wire \core_0.dec_rf_ie[4] ;
 wire \core_0.dec_rf_ie[5] ;
 wire \core_0.dec_rf_ie[6] ;
 wire \core_0.dec_rf_ie[7] ;
 wire \core_0.dec_sreg_irt ;
 wire \core_0.dec_sreg_jal_over ;
 wire \core_0.dec_sreg_load ;
 wire \core_0.dec_sreg_store ;
 wire \core_0.dec_sys ;
 wire \core_0.dec_used_operands[0] ;
 wire \core_0.dec_used_operands[1] ;
 wire \core_0.decode.i_flush ;
 wire \core_0.decode.i_imm_pass[0] ;
 wire \core_0.decode.i_imm_pass[10] ;
 wire \core_0.decode.i_imm_pass[11] ;
 wire \core_0.decode.i_imm_pass[12] ;
 wire \core_0.decode.i_imm_pass[13] ;
 wire \core_0.decode.i_imm_pass[14] ;
 wire \core_0.decode.i_imm_pass[15] ;
 wire \core_0.decode.i_imm_pass[1] ;
 wire \core_0.decode.i_imm_pass[2] ;
 wire \core_0.decode.i_imm_pass[3] ;
 wire \core_0.decode.i_imm_pass[4] ;
 wire \core_0.decode.i_imm_pass[5] ;
 wire \core_0.decode.i_imm_pass[6] ;
 wire \core_0.decode.i_imm_pass[7] ;
 wire \core_0.decode.i_imm_pass[8] ;
 wire \core_0.decode.i_imm_pass[9] ;
 wire \core_0.decode.i_instr_l[0] ;
 wire \core_0.decode.i_instr_l[10] ;
 wire \core_0.decode.i_instr_l[11] ;
 wire \core_0.decode.i_instr_l[12] ;
 wire \core_0.decode.i_instr_l[13] ;
 wire \core_0.decode.i_instr_l[14] ;
 wire \core_0.decode.i_instr_l[15] ;
 wire \core_0.decode.i_instr_l[1] ;
 wire \core_0.decode.i_instr_l[2] ;
 wire \core_0.decode.i_instr_l[3] ;
 wire \core_0.decode.i_instr_l[4] ;
 wire \core_0.decode.i_instr_l[5] ;
 wire \core_0.decode.i_instr_l[6] ;
 wire \core_0.decode.i_instr_l[7] ;
 wire \core_0.decode.i_instr_l[8] ;
 wire \core_0.decode.i_instr_l[9] ;
 wire \core_0.decode.i_jmp_pred_pass ;
 wire \core_0.decode.i_submit ;
 wire \core_0.decode.input_valid ;
 wire \core_0.decode.o_submit ;
 wire \core_0.decode.oc_alu_mode[11] ;
 wire \core_0.decode.oc_alu_mode[12] ;
 wire \core_0.decode.oc_alu_mode[13] ;
 wire \core_0.decode.oc_alu_mode[1] ;
 wire \core_0.decode.oc_alu_mode[2] ;
 wire \core_0.decode.oc_alu_mode[3] ;
 wire \core_0.decode.oc_alu_mode[4] ;
 wire \core_0.decode.oc_alu_mode[6] ;
 wire \core_0.decode.oc_alu_mode[7] ;
 wire \core_0.decode.oc_alu_mode[9] ;
 wire \core_0.ew_addr[0] ;
 wire \core_0.ew_addr_high[0] ;
 wire \core_0.ew_data[0] ;
 wire \core_0.ew_data[10] ;
 wire \core_0.ew_data[11] ;
 wire \core_0.ew_data[12] ;
 wire \core_0.ew_data[13] ;
 wire \core_0.ew_data[14] ;
 wire \core_0.ew_data[15] ;
 wire \core_0.ew_data[1] ;
 wire \core_0.ew_data[2] ;
 wire \core_0.ew_data[3] ;
 wire \core_0.ew_data[4] ;
 wire \core_0.ew_data[5] ;
 wire \core_0.ew_data[6] ;
 wire \core_0.ew_data[7] ;
 wire \core_0.ew_data[8] ;
 wire \core_0.ew_data[9] ;
 wire \core_0.ew_mem_access ;
 wire \core_0.ew_mem_width ;
 wire \core_0.ew_reg_ie[0] ;
 wire \core_0.ew_reg_ie[1] ;
 wire \core_0.ew_reg_ie[2] ;
 wire \core_0.ew_reg_ie[3] ;
 wire \core_0.ew_reg_ie[4] ;
 wire \core_0.ew_reg_ie[5] ;
 wire \core_0.ew_reg_ie[6] ;
 wire \core_0.ew_reg_ie[7] ;
 wire \core_0.ew_submit ;
 wire \core_0.execute.alu_flag_reg.o_d[0] ;
 wire \core_0.execute.alu_flag_reg.o_d[1] ;
 wire \core_0.execute.alu_flag_reg.o_d[2] ;
 wire \core_0.execute.alu_flag_reg.o_d[3] ;
 wire \core_0.execute.alu_flag_reg.o_d[4] ;
 wire \core_0.execute.alu_mul_div.cbit[0] ;
 wire \core_0.execute.alu_mul_div.cbit[1] ;
 wire \core_0.execute.alu_mul_div.cbit[2] ;
 wire \core_0.execute.alu_mul_div.cbit[3] ;
 wire \core_0.execute.alu_mul_div.comp ;
 wire \core_0.execute.alu_mul_div.div_cur[0] ;
 wire \core_0.execute.alu_mul_div.div_cur[10] ;
 wire \core_0.execute.alu_mul_div.div_cur[11] ;
 wire \core_0.execute.alu_mul_div.div_cur[12] ;
 wire \core_0.execute.alu_mul_div.div_cur[13] ;
 wire \core_0.execute.alu_mul_div.div_cur[14] ;
 wire \core_0.execute.alu_mul_div.div_cur[15] ;
 wire \core_0.execute.alu_mul_div.div_cur[1] ;
 wire \core_0.execute.alu_mul_div.div_cur[2] ;
 wire \core_0.execute.alu_mul_div.div_cur[3] ;
 wire \core_0.execute.alu_mul_div.div_cur[4] ;
 wire \core_0.execute.alu_mul_div.div_cur[5] ;
 wire \core_0.execute.alu_mul_div.div_cur[6] ;
 wire \core_0.execute.alu_mul_div.div_cur[7] ;
 wire \core_0.execute.alu_mul_div.div_cur[8] ;
 wire \core_0.execute.alu_mul_div.div_cur[9] ;
 wire \core_0.execute.alu_mul_div.div_res[0] ;
 wire \core_0.execute.alu_mul_div.div_res[10] ;
 wire \core_0.execute.alu_mul_div.div_res[11] ;
 wire \core_0.execute.alu_mul_div.div_res[12] ;
 wire \core_0.execute.alu_mul_div.div_res[13] ;
 wire \core_0.execute.alu_mul_div.div_res[14] ;
 wire \core_0.execute.alu_mul_div.div_res[15] ;
 wire \core_0.execute.alu_mul_div.div_res[1] ;
 wire \core_0.execute.alu_mul_div.div_res[2] ;
 wire \core_0.execute.alu_mul_div.div_res[3] ;
 wire \core_0.execute.alu_mul_div.div_res[4] ;
 wire \core_0.execute.alu_mul_div.div_res[5] ;
 wire \core_0.execute.alu_mul_div.div_res[6] ;
 wire \core_0.execute.alu_mul_div.div_res[7] ;
 wire \core_0.execute.alu_mul_div.div_res[8] ;
 wire \core_0.execute.alu_mul_div.div_res[9] ;
 wire \core_0.execute.alu_mul_div.i_div ;
 wire \core_0.execute.alu_mul_div.i_mod ;
 wire \core_0.execute.alu_mul_div.i_mul ;
 wire \core_0.execute.alu_mul_div.mul_res[0] ;
 wire \core_0.execute.alu_mul_div.mul_res[10] ;
 wire \core_0.execute.alu_mul_div.mul_res[11] ;
 wire \core_0.execute.alu_mul_div.mul_res[12] ;
 wire \core_0.execute.alu_mul_div.mul_res[13] ;
 wire \core_0.execute.alu_mul_div.mul_res[14] ;
 wire \core_0.execute.alu_mul_div.mul_res[15] ;
 wire \core_0.execute.alu_mul_div.mul_res[1] ;
 wire \core_0.execute.alu_mul_div.mul_res[2] ;
 wire \core_0.execute.alu_mul_div.mul_res[3] ;
 wire \core_0.execute.alu_mul_div.mul_res[4] ;
 wire \core_0.execute.alu_mul_div.mul_res[5] ;
 wire \core_0.execute.alu_mul_div.mul_res[6] ;
 wire \core_0.execute.alu_mul_div.mul_res[7] ;
 wire \core_0.execute.alu_mul_div.mul_res[8] ;
 wire \core_0.execute.alu_mul_div.mul_res[9] ;
 wire \core_0.execute.hold_valid ;
 wire \core_0.execute.irq_en ;
 wire \core_0.execute.mem_stage_pc[0] ;
 wire \core_0.execute.mem_stage_pc[10] ;
 wire \core_0.execute.mem_stage_pc[11] ;
 wire \core_0.execute.mem_stage_pc[12] ;
 wire \core_0.execute.mem_stage_pc[13] ;
 wire \core_0.execute.mem_stage_pc[14] ;
 wire \core_0.execute.mem_stage_pc[15] ;
 wire \core_0.execute.mem_stage_pc[1] ;
 wire \core_0.execute.mem_stage_pc[2] ;
 wire \core_0.execute.mem_stage_pc[3] ;
 wire \core_0.execute.mem_stage_pc[4] ;
 wire \core_0.execute.mem_stage_pc[5] ;
 wire \core_0.execute.mem_stage_pc[6] ;
 wire \core_0.execute.mem_stage_pc[7] ;
 wire \core_0.execute.mem_stage_pc[8] ;
 wire \core_0.execute.mem_stage_pc[9] ;
 wire \core_0.execute.next_ready_delayed ;
 wire \core_0.execute.pc_high_buff_out[0] ;
 wire \core_0.execute.pc_high_buff_out[1] ;
 wire \core_0.execute.pc_high_buff_out[2] ;
 wire \core_0.execute.pc_high_buff_out[3] ;
 wire \core_0.execute.pc_high_buff_out[4] ;
 wire \core_0.execute.pc_high_buff_out[5] ;
 wire \core_0.execute.pc_high_buff_out[6] ;
 wire \core_0.execute.pc_high_buff_out[7] ;
 wire \core_0.execute.pc_high_out[0] ;
 wire \core_0.execute.pc_high_out[1] ;
 wire \core_0.execute.pc_high_out[2] ;
 wire \core_0.execute.pc_high_out[3] ;
 wire \core_0.execute.pc_high_out[4] ;
 wire \core_0.execute.pc_high_out[5] ;
 wire \core_0.execute.pc_high_out[6] ;
 wire \core_0.execute.pc_high_out[7] ;
 wire \core_0.execute.prev_pc_high[0] ;
 wire \core_0.execute.prev_pc_high[1] ;
 wire \core_0.execute.prev_pc_high[2] ;
 wire \core_0.execute.prev_pc_high[3] ;
 wire \core_0.execute.prev_pc_high[4] ;
 wire \core_0.execute.prev_pc_high[5] ;
 wire \core_0.execute.prev_pc_high[6] ;
 wire \core_0.execute.prev_pc_high[7] ;
 wire \core_0.execute.prev_sys ;
 wire \core_0.execute.rf.reg_outputs[1][0] ;
 wire \core_0.execute.rf.reg_outputs[1][10] ;
 wire \core_0.execute.rf.reg_outputs[1][11] ;
 wire \core_0.execute.rf.reg_outputs[1][12] ;
 wire \core_0.execute.rf.reg_outputs[1][13] ;
 wire \core_0.execute.rf.reg_outputs[1][14] ;
 wire \core_0.execute.rf.reg_outputs[1][15] ;
 wire \core_0.execute.rf.reg_outputs[1][1] ;
 wire \core_0.execute.rf.reg_outputs[1][2] ;
 wire \core_0.execute.rf.reg_outputs[1][3] ;
 wire \core_0.execute.rf.reg_outputs[1][4] ;
 wire \core_0.execute.rf.reg_outputs[1][5] ;
 wire \core_0.execute.rf.reg_outputs[1][6] ;
 wire \core_0.execute.rf.reg_outputs[1][7] ;
 wire \core_0.execute.rf.reg_outputs[1][8] ;
 wire \core_0.execute.rf.reg_outputs[1][9] ;
 wire \core_0.execute.rf.reg_outputs[2][0] ;
 wire \core_0.execute.rf.reg_outputs[2][10] ;
 wire \core_0.execute.rf.reg_outputs[2][11] ;
 wire \core_0.execute.rf.reg_outputs[2][12] ;
 wire \core_0.execute.rf.reg_outputs[2][13] ;
 wire \core_0.execute.rf.reg_outputs[2][14] ;
 wire \core_0.execute.rf.reg_outputs[2][15] ;
 wire \core_0.execute.rf.reg_outputs[2][1] ;
 wire \core_0.execute.rf.reg_outputs[2][2] ;
 wire \core_0.execute.rf.reg_outputs[2][3] ;
 wire \core_0.execute.rf.reg_outputs[2][4] ;
 wire \core_0.execute.rf.reg_outputs[2][5] ;
 wire \core_0.execute.rf.reg_outputs[2][6] ;
 wire \core_0.execute.rf.reg_outputs[2][7] ;
 wire \core_0.execute.rf.reg_outputs[2][8] ;
 wire \core_0.execute.rf.reg_outputs[2][9] ;
 wire \core_0.execute.rf.reg_outputs[3][0] ;
 wire \core_0.execute.rf.reg_outputs[3][10] ;
 wire \core_0.execute.rf.reg_outputs[3][11] ;
 wire \core_0.execute.rf.reg_outputs[3][12] ;
 wire \core_0.execute.rf.reg_outputs[3][13] ;
 wire \core_0.execute.rf.reg_outputs[3][14] ;
 wire \core_0.execute.rf.reg_outputs[3][15] ;
 wire \core_0.execute.rf.reg_outputs[3][1] ;
 wire \core_0.execute.rf.reg_outputs[3][2] ;
 wire \core_0.execute.rf.reg_outputs[3][3] ;
 wire \core_0.execute.rf.reg_outputs[3][4] ;
 wire \core_0.execute.rf.reg_outputs[3][5] ;
 wire \core_0.execute.rf.reg_outputs[3][6] ;
 wire \core_0.execute.rf.reg_outputs[3][7] ;
 wire \core_0.execute.rf.reg_outputs[3][8] ;
 wire \core_0.execute.rf.reg_outputs[3][9] ;
 wire \core_0.execute.rf.reg_outputs[4][0] ;
 wire \core_0.execute.rf.reg_outputs[4][10] ;
 wire \core_0.execute.rf.reg_outputs[4][11] ;
 wire \core_0.execute.rf.reg_outputs[4][12] ;
 wire \core_0.execute.rf.reg_outputs[4][13] ;
 wire \core_0.execute.rf.reg_outputs[4][14] ;
 wire \core_0.execute.rf.reg_outputs[4][15] ;
 wire \core_0.execute.rf.reg_outputs[4][1] ;
 wire \core_0.execute.rf.reg_outputs[4][2] ;
 wire \core_0.execute.rf.reg_outputs[4][3] ;
 wire \core_0.execute.rf.reg_outputs[4][4] ;
 wire \core_0.execute.rf.reg_outputs[4][5] ;
 wire \core_0.execute.rf.reg_outputs[4][6] ;
 wire \core_0.execute.rf.reg_outputs[4][7] ;
 wire \core_0.execute.rf.reg_outputs[4][8] ;
 wire \core_0.execute.rf.reg_outputs[4][9] ;
 wire \core_0.execute.rf.reg_outputs[5][0] ;
 wire \core_0.execute.rf.reg_outputs[5][10] ;
 wire \core_0.execute.rf.reg_outputs[5][11] ;
 wire \core_0.execute.rf.reg_outputs[5][12] ;
 wire \core_0.execute.rf.reg_outputs[5][13] ;
 wire \core_0.execute.rf.reg_outputs[5][14] ;
 wire \core_0.execute.rf.reg_outputs[5][15] ;
 wire \core_0.execute.rf.reg_outputs[5][1] ;
 wire \core_0.execute.rf.reg_outputs[5][2] ;
 wire \core_0.execute.rf.reg_outputs[5][3] ;
 wire \core_0.execute.rf.reg_outputs[5][4] ;
 wire \core_0.execute.rf.reg_outputs[5][5] ;
 wire \core_0.execute.rf.reg_outputs[5][6] ;
 wire \core_0.execute.rf.reg_outputs[5][7] ;
 wire \core_0.execute.rf.reg_outputs[5][8] ;
 wire \core_0.execute.rf.reg_outputs[5][9] ;
 wire \core_0.execute.rf.reg_outputs[6][0] ;
 wire \core_0.execute.rf.reg_outputs[6][10] ;
 wire \core_0.execute.rf.reg_outputs[6][11] ;
 wire \core_0.execute.rf.reg_outputs[6][12] ;
 wire \core_0.execute.rf.reg_outputs[6][13] ;
 wire \core_0.execute.rf.reg_outputs[6][14] ;
 wire \core_0.execute.rf.reg_outputs[6][15] ;
 wire \core_0.execute.rf.reg_outputs[6][1] ;
 wire \core_0.execute.rf.reg_outputs[6][2] ;
 wire \core_0.execute.rf.reg_outputs[6][3] ;
 wire \core_0.execute.rf.reg_outputs[6][4] ;
 wire \core_0.execute.rf.reg_outputs[6][5] ;
 wire \core_0.execute.rf.reg_outputs[6][6] ;
 wire \core_0.execute.rf.reg_outputs[6][7] ;
 wire \core_0.execute.rf.reg_outputs[6][8] ;
 wire \core_0.execute.rf.reg_outputs[6][9] ;
 wire \core_0.execute.rf.reg_outputs[7][0] ;
 wire \core_0.execute.rf.reg_outputs[7][10] ;
 wire \core_0.execute.rf.reg_outputs[7][11] ;
 wire \core_0.execute.rf.reg_outputs[7][12] ;
 wire \core_0.execute.rf.reg_outputs[7][13] ;
 wire \core_0.execute.rf.reg_outputs[7][14] ;
 wire \core_0.execute.rf.reg_outputs[7][15] ;
 wire \core_0.execute.rf.reg_outputs[7][1] ;
 wire \core_0.execute.rf.reg_outputs[7][2] ;
 wire \core_0.execute.rf.reg_outputs[7][3] ;
 wire \core_0.execute.rf.reg_outputs[7][4] ;
 wire \core_0.execute.rf.reg_outputs[7][5] ;
 wire \core_0.execute.rf.reg_outputs[7][6] ;
 wire \core_0.execute.rf.reg_outputs[7][7] ;
 wire \core_0.execute.rf.reg_outputs[7][8] ;
 wire \core_0.execute.rf.reg_outputs[7][9] ;
 wire \core_0.execute.sreg_data_page ;
 wire \core_0.execute.sreg_irq_flags.i_d[2] ;
 wire \core_0.execute.sreg_irq_flags.o_d[0] ;
 wire \core_0.execute.sreg_irq_flags.o_d[1] ;
 wire \core_0.execute.sreg_irq_flags.o_d[2] ;
 wire \core_0.execute.sreg_irq_flags.o_d[3] ;
 wire \core_0.execute.sreg_irq_flags.o_d[4] ;
 wire \core_0.execute.sreg_irq_pc.o_d[0] ;
 wire \core_0.execute.sreg_irq_pc.o_d[10] ;
 wire \core_0.execute.sreg_irq_pc.o_d[11] ;
 wire \core_0.execute.sreg_irq_pc.o_d[12] ;
 wire \core_0.execute.sreg_irq_pc.o_d[13] ;
 wire \core_0.execute.sreg_irq_pc.o_d[14] ;
 wire \core_0.execute.sreg_irq_pc.o_d[15] ;
 wire \core_0.execute.sreg_irq_pc.o_d[1] ;
 wire \core_0.execute.sreg_irq_pc.o_d[2] ;
 wire \core_0.execute.sreg_irq_pc.o_d[3] ;
 wire \core_0.execute.sreg_irq_pc.o_d[4] ;
 wire \core_0.execute.sreg_irq_pc.o_d[5] ;
 wire \core_0.execute.sreg_irq_pc.o_d[6] ;
 wire \core_0.execute.sreg_irq_pc.o_d[7] ;
 wire \core_0.execute.sreg_irq_pc.o_d[8] ;
 wire \core_0.execute.sreg_irq_pc.o_d[9] ;
 wire \core_0.execute.sreg_jtr_buff.o_d[0] ;
 wire \core_0.execute.sreg_jtr_buff.o_d[1] ;
 wire \core_0.execute.sreg_jtr_buff.o_d[2] ;
 wire \core_0.execute.sreg_long_ptr_en ;
 wire \core_0.execute.sreg_priv_control.o_d[0] ;
 wire \core_0.execute.sreg_priv_control.o_d[10] ;
 wire \core_0.execute.sreg_priv_control.o_d[11] ;
 wire \core_0.execute.sreg_priv_control.o_d[12] ;
 wire \core_0.execute.sreg_priv_control.o_d[13] ;
 wire \core_0.execute.sreg_priv_control.o_d[14] ;
 wire \core_0.execute.sreg_priv_control.o_d[15] ;
 wire \core_0.execute.sreg_priv_control.o_d[4] ;
 wire \core_0.execute.sreg_priv_control.o_d[5] ;
 wire \core_0.execute.sreg_priv_control.o_d[6] ;
 wire \core_0.execute.sreg_priv_control.o_d[7] ;
 wire \core_0.execute.sreg_priv_control.o_d[8] ;
 wire \core_0.execute.sreg_priv_control.o_d[9] ;
 wire \core_0.execute.sreg_scratch.o_d[0] ;
 wire \core_0.execute.sreg_scratch.o_d[10] ;
 wire \core_0.execute.sreg_scratch.o_d[11] ;
 wire \core_0.execute.sreg_scratch.o_d[12] ;
 wire \core_0.execute.sreg_scratch.o_d[13] ;
 wire \core_0.execute.sreg_scratch.o_d[14] ;
 wire \core_0.execute.sreg_scratch.o_d[15] ;
 wire \core_0.execute.sreg_scratch.o_d[1] ;
 wire \core_0.execute.sreg_scratch.o_d[2] ;
 wire \core_0.execute.sreg_scratch.o_d[3] ;
 wire \core_0.execute.sreg_scratch.o_d[4] ;
 wire \core_0.execute.sreg_scratch.o_d[5] ;
 wire \core_0.execute.sreg_scratch.o_d[6] ;
 wire \core_0.execute.sreg_scratch.o_d[7] ;
 wire \core_0.execute.sreg_scratch.o_d[8] ;
 wire \core_0.execute.sreg_scratch.o_d[9] ;
 wire \core_0.execute.trap_flag ;
 wire \core_0.fetch.current_req_branch_pred ;
 wire \core_0.fetch.dbg_out ;
 wire \core_0.fetch.flush_event_invalidate ;
 wire \core_0.fetch.out_buffer_data_instr[0] ;
 wire \core_0.fetch.out_buffer_data_instr[10] ;
 wire \core_0.fetch.out_buffer_data_instr[11] ;
 wire \core_0.fetch.out_buffer_data_instr[12] ;
 wire \core_0.fetch.out_buffer_data_instr[13] ;
 wire \core_0.fetch.out_buffer_data_instr[14] ;
 wire \core_0.fetch.out_buffer_data_instr[15] ;
 wire \core_0.fetch.out_buffer_data_instr[16] ;
 wire \core_0.fetch.out_buffer_data_instr[17] ;
 wire \core_0.fetch.out_buffer_data_instr[18] ;
 wire \core_0.fetch.out_buffer_data_instr[19] ;
 wire \core_0.fetch.out_buffer_data_instr[1] ;
 wire \core_0.fetch.out_buffer_data_instr[20] ;
 wire \core_0.fetch.out_buffer_data_instr[21] ;
 wire \core_0.fetch.out_buffer_data_instr[22] ;
 wire \core_0.fetch.out_buffer_data_instr[23] ;
 wire \core_0.fetch.out_buffer_data_instr[24] ;
 wire \core_0.fetch.out_buffer_data_instr[25] ;
 wire \core_0.fetch.out_buffer_data_instr[26] ;
 wire \core_0.fetch.out_buffer_data_instr[27] ;
 wire \core_0.fetch.out_buffer_data_instr[28] ;
 wire \core_0.fetch.out_buffer_data_instr[29] ;
 wire \core_0.fetch.out_buffer_data_instr[2] ;
 wire \core_0.fetch.out_buffer_data_instr[30] ;
 wire \core_0.fetch.out_buffer_data_instr[31] ;
 wire \core_0.fetch.out_buffer_data_instr[3] ;
 wire \core_0.fetch.out_buffer_data_instr[4] ;
 wire \core_0.fetch.out_buffer_data_instr[5] ;
 wire \core_0.fetch.out_buffer_data_instr[6] ;
 wire \core_0.fetch.out_buffer_data_instr[7] ;
 wire \core_0.fetch.out_buffer_data_instr[8] ;
 wire \core_0.fetch.out_buffer_data_instr[9] ;
 wire \core_0.fetch.out_buffer_data_pred ;
 wire \core_0.fetch.out_buffer_valid ;
 wire \core_0.fetch.pc_flush_override ;
 wire \core_0.fetch.pc_reset_override ;
 wire \core_0.fetch.prev_req_branch_pred ;
 wire \core_0.fetch.prev_request_pc[0] ;
 wire \core_0.fetch.prev_request_pc[10] ;
 wire \core_0.fetch.prev_request_pc[11] ;
 wire \core_0.fetch.prev_request_pc[12] ;
 wire \core_0.fetch.prev_request_pc[13] ;
 wire \core_0.fetch.prev_request_pc[14] ;
 wire \core_0.fetch.prev_request_pc[15] ;
 wire \core_0.fetch.prev_request_pc[1] ;
 wire \core_0.fetch.prev_request_pc[2] ;
 wire \core_0.fetch.prev_request_pc[3] ;
 wire \core_0.fetch.prev_request_pc[4] ;
 wire \core_0.fetch.prev_request_pc[5] ;
 wire \core_0.fetch.prev_request_pc[6] ;
 wire \core_0.fetch.prev_request_pc[7] ;
 wire \core_0.fetch.prev_request_pc[8] ;
 wire \core_0.fetch.prev_request_pc[9] ;
 wire \core_0.fetch.submitable ;
 wire clknet_leaf_0_i_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_9_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_0_i_clk;
 wire clknet_1_0_0_i_clk;
 wire clknet_1_0_1_i_clk;
 wire clknet_1_1_0_i_clk;
 wire clknet_1_1_1_i_clk;
 wire clknet_2_0_0_i_clk;
 wire clknet_2_1_0_i_clk;
 wire clknet_2_2_0_i_clk;
 wire clknet_2_3_0_i_clk;
 wire clknet_opt_1_0_i_clk;
 wire clknet_opt_1_1_i_clk;

 sky130_fd_sc_hd__buf_2 _3408_ (.A(\core_0.dec_r_reg_sel[2] ),
    .X(_0515_));
 sky130_fd_sc_hd__clkbuf_2 _3409_ (.A(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_2 _3410_ (.A(\core_0.dec_r_reg_sel[1] ),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_2 _3411_ (.A(\core_0.dec_r_reg_sel[0] ),
    .X(_0518_));
 sky130_fd_sc_hd__or3_1 _3412_ (.A(_0516_),
    .B(_0517_),
    .C(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__buf_6 _3413_ (.A(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__buf_6 _3414_ (.A(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__and3b_1 _3415_ (.A_N(_0516_),
    .B(_0517_),
    .C(_0518_),
    .X(_0522_));
 sky130_fd_sc_hd__buf_2 _3416_ (.A(\core_0.dec_r_reg_sel[2] ),
    .X(_0523_));
 sky130_fd_sc_hd__buf_2 _3417_ (.A(\core_0.dec_r_reg_sel[0] ),
    .X(_0524_));
 sky130_fd_sc_hd__nor3b_4 _3418_ (.A(_0523_),
    .B(_0524_),
    .C_N(\core_0.dec_r_reg_sel[1] ),
    .Y(_0525_));
 sky130_fd_sc_hd__buf_4 _3419_ (.A(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__buf_2 _3420_ (.A(\core_0.dec_r_reg_sel[0] ),
    .X(_0527_));
 sky130_fd_sc_hd__and4_1 _3421_ (.A(\core_0.execute.rf.reg_outputs[7][15] ),
    .B(_0516_),
    .C(_0517_),
    .D(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__a221o_1 _3422_ (.A1(\core_0.execute.rf.reg_outputs[3][15] ),
    .A2(_0522_),
    .B1(_0526_),
    .B2(\core_0.execute.rf.reg_outputs[2][15] ),
    .C1(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__buf_2 _3423_ (.A(_0517_),
    .X(_0530_));
 sky130_fd_sc_hd__buf_2 _3424_ (.A(_0518_),
    .X(_0531_));
 sky130_fd_sc_hd__nor2_1 _3425_ (.A(_0530_),
    .B(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__or2b_1 _3426_ (.A(\core_0.execute.rf.reg_outputs[4][15] ),
    .B_N(_0516_),
    .X(_0533_));
 sky130_fd_sc_hd__and4b_1 _3427_ (.A_N(_0517_),
    .B(_0518_),
    .C(\core_0.execute.rf.reg_outputs[5][15] ),
    .D(_0516_),
    .X(_0534_));
 sky130_fd_sc_hd__and4b_1 _3428_ (.A_N(_0518_),
    .B(_0517_),
    .C(_0516_),
    .D(\core_0.execute.rf.reg_outputs[6][15] ),
    .X(_0535_));
 sky130_fd_sc_hd__buf_2 _3429_ (.A(_0515_),
    .X(_0536_));
 sky130_fd_sc_hd__buf_2 _3430_ (.A(\core_0.dec_r_reg_sel[1] ),
    .X(_0537_));
 sky130_fd_sc_hd__clkbuf_2 _3431_ (.A(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__and4bb_1 _3432_ (.A_N(_0536_),
    .B_N(_0538_),
    .C(_0518_),
    .D(\core_0.execute.rf.reg_outputs[1][15] ),
    .X(_0539_));
 sky130_fd_sc_hd__a2111o_1 _3433_ (.A1(_0532_),
    .A2(_0533_),
    .B1(_0534_),
    .C1(_0535_),
    .D1(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__o22a_1 _3434_ (.A1(net94),
    .A2(_0521_),
    .B1(_0529_),
    .B2(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__buf_6 _3435_ (.A(_0541_),
    .X(net200));
 sky130_fd_sc_hd__nor3b_4 _3436_ (.A(_0515_),
    .B(_0537_),
    .C_N(\core_0.dec_r_reg_sel[0] ),
    .Y(_0542_));
 sky130_fd_sc_hd__and4b_1 _3437_ (.A_N(_0527_),
    .B(_0538_),
    .C(_0536_),
    .D(\core_0.execute.rf.reg_outputs[6][14] ),
    .X(_0543_));
 sky130_fd_sc_hd__a221o_1 _3438_ (.A1(\core_0.execute.rf.reg_outputs[3][14] ),
    .A2(_0522_),
    .B1(_0542_),
    .B2(\core_0.execute.rf.reg_outputs[1][14] ),
    .C1(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__and3_1 _3439_ (.A(_0536_),
    .B(_0517_),
    .C(_0527_),
    .X(_0545_));
 sky130_fd_sc_hd__buf_2 _3440_ (.A(_0516_),
    .X(_0546_));
 sky130_fd_sc_hd__or2b_1 _3441_ (.A(\core_0.execute.rf.reg_outputs[4][14] ),
    .B_N(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__a22o_1 _3442_ (.A1(\core_0.execute.rf.reg_outputs[7][14] ),
    .A2(_0545_),
    .B1(_0547_),
    .B2(_0532_),
    .X(_0548_));
 sky130_fd_sc_hd__and3b_1 _3443_ (.A_N(\core_0.dec_r_reg_sel[1] ),
    .B(\core_0.dec_r_reg_sel[0] ),
    .C(_0515_),
    .X(_0549_));
 sky130_fd_sc_hd__clkbuf_4 _3444_ (.A(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__a22o_1 _3445_ (.A1(\core_0.execute.rf.reg_outputs[2][14] ),
    .A2(_0526_),
    .B1(_0550_),
    .B2(\core_0.execute.rf.reg_outputs[5][14] ),
    .X(_0551_));
 sky130_fd_sc_hd__or2_1 _3446_ (.A(net93),
    .B(_0519_),
    .X(_0552_));
 sky130_fd_sc_hd__o31a_1 _3447_ (.A1(_0544_),
    .A2(_0548_),
    .A3(_0551_),
    .B1(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__buf_6 _3448_ (.A(_0553_),
    .X(net199));
 sky130_fd_sc_hd__nor3b_1 _3449_ (.A(\core_0.dec_r_reg_sel[1] ),
    .B(\core_0.dec_r_reg_sel[0] ),
    .C_N(_0515_),
    .Y(_0554_));
 sky130_fd_sc_hd__buf_4 _3450_ (.A(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__buf_2 _3451_ (.A(_0523_),
    .X(_0556_));
 sky130_fd_sc_hd__buf_2 _3452_ (.A(_0517_),
    .X(_0557_));
 sky130_fd_sc_hd__buf_2 _3453_ (.A(_0524_),
    .X(_0558_));
 sky130_fd_sc_hd__and4bb_1 _3454_ (.A_N(_0556_),
    .B_N(_0557_),
    .C(_0558_),
    .D(\core_0.execute.rf.reg_outputs[1][13] ),
    .X(_0559_));
 sky130_fd_sc_hd__and4b_1 _3455_ (.A_N(_0530_),
    .B(_0558_),
    .C(\core_0.execute.rf.reg_outputs[5][13] ),
    .D(_0556_),
    .X(_0560_));
 sky130_fd_sc_hd__and4b_1 _3456_ (.A_N(_0531_),
    .B(_0530_),
    .C(_0546_),
    .D(\core_0.execute.rf.reg_outputs[6][13] ),
    .X(_0561_));
 sky130_fd_sc_hd__a2111o_1 _3457_ (.A1(\core_0.execute.rf.reg_outputs[4][13] ),
    .A2(_0555_),
    .B1(_0559_),
    .C1(_0560_),
    .D1(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__and4b_1 _3458_ (.A_N(_0556_),
    .B(_0557_),
    .C(_0558_),
    .D(\core_0.execute.rf.reg_outputs[3][13] ),
    .X(_0563_));
 sky130_fd_sc_hd__and4_1 _3459_ (.A(\core_0.execute.rf.reg_outputs[7][13] ),
    .B(_0556_),
    .C(_0557_),
    .D(_0558_),
    .X(_0564_));
 sky130_fd_sc_hd__nor3_2 _3460_ (.A(_0515_),
    .B(\core_0.dec_r_reg_sel[1] ),
    .C(\core_0.dec_r_reg_sel[0] ),
    .Y(_0565_));
 sky130_fd_sc_hd__buf_4 _3461_ (.A(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__a2111o_1 _3462_ (.A1(\core_0.execute.rf.reg_outputs[2][13] ),
    .A2(_0526_),
    .B1(_0563_),
    .C1(_0564_),
    .D1(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__o22a_1 _3463_ (.A1(net92),
    .A2(_0521_),
    .B1(_0562_),
    .B2(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__buf_6 _3464_ (.A(_0568_),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 _3465_ (.A(_0537_),
    .X(_0569_));
 sky130_fd_sc_hd__and4b_1 _3466_ (.A_N(_0569_),
    .B(_0531_),
    .C(\core_0.execute.rf.reg_outputs[5][12] ),
    .D(_0546_),
    .X(_0570_));
 sky130_fd_sc_hd__clkbuf_4 _3467_ (.A(_0518_),
    .X(_0571_));
 sky130_fd_sc_hd__and4b_1 _3468_ (.A_N(_0571_),
    .B(_0530_),
    .C(_0546_),
    .D(\core_0.execute.rf.reg_outputs[6][12] ),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_4 _3469_ (.A(_0523_),
    .X(_0573_));
 sky130_fd_sc_hd__and4bb_1 _3470_ (.A_N(_0573_),
    .B_N(_0569_),
    .C(_0571_),
    .D(\core_0.execute.rf.reg_outputs[1][12] ),
    .X(_0574_));
 sky130_fd_sc_hd__a2111o_2 _3471_ (.A1(\core_0.execute.rf.reg_outputs[4][12] ),
    .A2(_0555_),
    .B1(_0570_),
    .C1(_0572_),
    .D1(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__and4_1 _3472_ (.A(\core_0.execute.rf.reg_outputs[7][12] ),
    .B(_0546_),
    .C(_0530_),
    .D(_0531_),
    .X(_0576_));
 sky130_fd_sc_hd__and4b_1 _3473_ (.A_N(_0573_),
    .B(_0530_),
    .C(_0531_),
    .D(\core_0.execute.rf.reg_outputs[3][12] ),
    .X(_0577_));
 sky130_fd_sc_hd__a2111o_2 _3474_ (.A1(\core_0.execute.rf.reg_outputs[2][12] ),
    .A2(_0526_),
    .B1(_0576_),
    .C1(_0577_),
    .D1(_0566_),
    .X(_0578_));
 sky130_fd_sc_hd__o22ai_4 _3475_ (.A1(net91),
    .A2(_0521_),
    .B1(_0575_),
    .B2(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__clkinv_4 _3476_ (.A(_0579_),
    .Y(net197));
 sky130_fd_sc_hd__a22o_1 _3477_ (.A1(\core_0.execute.rf.reg_outputs[5][11] ),
    .A2(_0550_),
    .B1(_0555_),
    .B2(\core_0.execute.rf.reg_outputs[4][11] ),
    .X(_0580_));
 sky130_fd_sc_hd__and3b_4 _3478_ (.A_N(_0524_),
    .B(_0537_),
    .C(_0523_),
    .X(_0581_));
 sky130_fd_sc_hd__a22o_1 _3479_ (.A1(\core_0.execute.rf.reg_outputs[1][11] ),
    .A2(_0542_),
    .B1(_0581_),
    .B2(\core_0.execute.rf.reg_outputs[6][11] ),
    .X(_0582_));
 sky130_fd_sc_hd__and4b_1 _3480_ (.A_N(_0523_),
    .B(_0537_),
    .C(_0524_),
    .D(\core_0.execute.rf.reg_outputs[3][11] ),
    .X(_0583_));
 sky130_fd_sc_hd__and4_1 _3481_ (.A(\core_0.execute.rf.reg_outputs[7][11] ),
    .B(_0523_),
    .C(_0537_),
    .D(_0524_),
    .X(_0584_));
 sky130_fd_sc_hd__a2111o_1 _3482_ (.A1(\core_0.execute.rf.reg_outputs[2][11] ),
    .A2(_0525_),
    .B1(_0583_),
    .C1(_0584_),
    .D1(_0565_),
    .X(_0585_));
 sky130_fd_sc_hd__o32a_1 _3483_ (.A1(_0580_),
    .A2(_0582_),
    .A3(_0585_),
    .B1(_0520_),
    .B2(net90),
    .X(_0586_));
 sky130_fd_sc_hd__clkbuf_8 _3484_ (.A(_0586_),
    .X(net196));
 sky130_fd_sc_hd__a22o_1 _3485_ (.A1(\core_0.execute.rf.reg_outputs[5][10] ),
    .A2(_0550_),
    .B1(_0554_),
    .B2(\core_0.execute.rf.reg_outputs[4][10] ),
    .X(_0587_));
 sky130_fd_sc_hd__a22o_1 _3486_ (.A1(\core_0.execute.rf.reg_outputs[1][10] ),
    .A2(_0542_),
    .B1(_0581_),
    .B2(\core_0.execute.rf.reg_outputs[6][10] ),
    .X(_0588_));
 sky130_fd_sc_hd__and4b_1 _3487_ (.A_N(_0515_),
    .B(\core_0.dec_r_reg_sel[1] ),
    .C(\core_0.dec_r_reg_sel[0] ),
    .D(\core_0.execute.rf.reg_outputs[3][10] ),
    .X(_0589_));
 sky130_fd_sc_hd__and4_1 _3488_ (.A(\core_0.execute.rf.reg_outputs[7][10] ),
    .B(_0515_),
    .C(\core_0.dec_r_reg_sel[1] ),
    .D(_0524_),
    .X(_0590_));
 sky130_fd_sc_hd__a2111o_1 _3489_ (.A1(\core_0.execute.rf.reg_outputs[2][10] ),
    .A2(_0525_),
    .B1(_0589_),
    .C1(_0590_),
    .D1(_0565_),
    .X(_0591_));
 sky130_fd_sc_hd__o32ai_4 _3490_ (.A1(_0587_),
    .A2(_0588_),
    .A3(_0591_),
    .B1(_0520_),
    .B2(net89),
    .Y(_0592_));
 sky130_fd_sc_hd__clkinv_4 _3491_ (.A(_0592_),
    .Y(net195));
 sky130_fd_sc_hd__a22o_1 _3492_ (.A1(\core_0.execute.rf.reg_outputs[5][9] ),
    .A2(_0550_),
    .B1(_0554_),
    .B2(\core_0.execute.rf.reg_outputs[4][9] ),
    .X(_0593_));
 sky130_fd_sc_hd__a22o_1 _3493_ (.A1(\core_0.execute.rf.reg_outputs[1][9] ),
    .A2(_0542_),
    .B1(_0581_),
    .B2(\core_0.execute.rf.reg_outputs[6][9] ),
    .X(_0594_));
 sky130_fd_sc_hd__and4b_1 _3494_ (.A_N(_0515_),
    .B(\core_0.dec_r_reg_sel[1] ),
    .C(\core_0.dec_r_reg_sel[0] ),
    .D(\core_0.execute.rf.reg_outputs[3][9] ),
    .X(_0595_));
 sky130_fd_sc_hd__and4_1 _3495_ (.A(\core_0.execute.rf.reg_outputs[7][9] ),
    .B(_0515_),
    .C(_0537_),
    .D(_0524_),
    .X(_0596_));
 sky130_fd_sc_hd__a2111o_1 _3496_ (.A1(\core_0.execute.rf.reg_outputs[2][9] ),
    .A2(_0525_),
    .B1(_0595_),
    .C1(_0596_),
    .D1(_0565_),
    .X(_0597_));
 sky130_fd_sc_hd__o32ai_4 _3497_ (.A1(_0593_),
    .A2(_0594_),
    .A3(_0597_),
    .B1(_0520_),
    .B2(net103),
    .Y(_0598_));
 sky130_fd_sc_hd__inv_4 _3498_ (.A(_0598_),
    .Y(net209));
 sky130_fd_sc_hd__a22o_1 _3499_ (.A1(\core_0.execute.rf.reg_outputs[5][8] ),
    .A2(_0550_),
    .B1(_0555_),
    .B2(\core_0.execute.rf.reg_outputs[4][8] ),
    .X(_0599_));
 sky130_fd_sc_hd__a22o_1 _3500_ (.A1(\core_0.execute.rf.reg_outputs[1][8] ),
    .A2(_0542_),
    .B1(_0581_),
    .B2(\core_0.execute.rf.reg_outputs[6][8] ),
    .X(_0600_));
 sky130_fd_sc_hd__and4b_1 _3501_ (.A_N(_0523_),
    .B(_0537_),
    .C(_0524_),
    .D(\core_0.execute.rf.reg_outputs[3][8] ),
    .X(_0601_));
 sky130_fd_sc_hd__and4_1 _3502_ (.A(\core_0.execute.rf.reg_outputs[7][8] ),
    .B(_0523_),
    .C(_0537_),
    .D(_0524_),
    .X(_0602_));
 sky130_fd_sc_hd__a2111o_1 _3503_ (.A1(\core_0.execute.rf.reg_outputs[2][8] ),
    .A2(_0525_),
    .B1(_0601_),
    .C1(_0602_),
    .D1(_0566_),
    .X(_0603_));
 sky130_fd_sc_hd__o32ai_4 _3504_ (.A1(_0599_),
    .A2(_0600_),
    .A3(_0603_),
    .B1(_0520_),
    .B2(net102),
    .Y(_0604_));
 sky130_fd_sc_hd__inv_4 _3505_ (.A(_0604_),
    .Y(net208));
 sky130_fd_sc_hd__and4_1 _3506_ (.A(\core_0.execute.rf.reg_outputs[7][7] ),
    .B(_0536_),
    .C(_0538_),
    .D(_0527_),
    .X(_0605_));
 sky130_fd_sc_hd__and4b_1 _3507_ (.A_N(_0556_),
    .B(_0538_),
    .C(_0527_),
    .D(\core_0.execute.rf.reg_outputs[3][7] ),
    .X(_0606_));
 sky130_fd_sc_hd__and4bb_1 _3508_ (.A_N(_0556_),
    .B_N(_0557_),
    .C(_0558_),
    .D(\core_0.execute.rf.reg_outputs[1][7] ),
    .X(_0607_));
 sky130_fd_sc_hd__a2111o_2 _3509_ (.A1(\core_0.execute.rf.reg_outputs[5][7] ),
    .A2(_0550_),
    .B1(_0605_),
    .C1(_0606_),
    .D1(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__and4bb_1 _3510_ (.A_N(_0538_),
    .B_N(_0527_),
    .C(\core_0.execute.rf.reg_outputs[4][7] ),
    .D(_0536_),
    .X(_0609_));
 sky130_fd_sc_hd__and4b_1 _3511_ (.A_N(_0558_),
    .B(_0538_),
    .C(_0536_),
    .D(\core_0.execute.rf.reg_outputs[6][7] ),
    .X(_0610_));
 sky130_fd_sc_hd__a2111o_2 _3512_ (.A1(\core_0.execute.rf.reg_outputs[2][7] ),
    .A2(_0526_),
    .B1(_0609_),
    .C1(_0610_),
    .D1(_0566_),
    .X(_0611_));
 sky130_fd_sc_hd__or2_1 _3513_ (.A(net101),
    .B(_0520_),
    .X(_0612_));
 sky130_fd_sc_hd__o21ai_4 _3514_ (.A1(_0608_),
    .A2(_0611_),
    .B1(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__inv_6 _3515_ (.A(_0613_),
    .Y(net207));
 sky130_fd_sc_hd__and4b_1 _3516_ (.A_N(_0557_),
    .B(_0527_),
    .C(\core_0.execute.rf.reg_outputs[5][6] ),
    .D(_0536_),
    .X(_0614_));
 sky130_fd_sc_hd__and4b_1 _3517_ (.A_N(_0531_),
    .B(_0557_),
    .C(_0556_),
    .D(\core_0.execute.rf.reg_outputs[6][6] ),
    .X(_0615_));
 sky130_fd_sc_hd__and4_1 _3518_ (.A(\core_0.execute.rf.reg_outputs[7][6] ),
    .B(_0556_),
    .C(_0530_),
    .D(_0531_),
    .X(_0616_));
 sky130_fd_sc_hd__a2111o_1 _3519_ (.A1(\core_0.execute.rf.reg_outputs[4][6] ),
    .A2(_0555_),
    .B1(_0614_),
    .C1(_0615_),
    .D1(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__a22o_1 _3520_ (.A1(\core_0.execute.rf.reg_outputs[2][6] ),
    .A2(_0526_),
    .B1(_0542_),
    .B2(\core_0.execute.rf.reg_outputs[1][6] ),
    .X(_0618_));
 sky130_fd_sc_hd__a21o_1 _3521_ (.A1(\core_0.execute.rf.reg_outputs[3][6] ),
    .A2(_0522_),
    .B1(_0566_),
    .X(_0619_));
 sky130_fd_sc_hd__or2_1 _3522_ (.A(net100),
    .B(_0520_),
    .X(_0620_));
 sky130_fd_sc_hd__o31a_1 _3523_ (.A1(_0617_),
    .A2(_0618_),
    .A3(_0619_),
    .B1(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__buf_8 _3524_ (.A(_0621_),
    .X(net206));
 sky130_fd_sc_hd__a22o_1 _3525_ (.A1(\core_0.execute.rf.reg_outputs[5][5] ),
    .A2(_0550_),
    .B1(_0555_),
    .B2(\core_0.execute.rf.reg_outputs[4][5] ),
    .X(_0622_));
 sky130_fd_sc_hd__a22o_1 _3526_ (.A1(\core_0.execute.rf.reg_outputs[1][5] ),
    .A2(_0542_),
    .B1(_0581_),
    .B2(\core_0.execute.rf.reg_outputs[6][5] ),
    .X(_0623_));
 sky130_fd_sc_hd__and4b_1 _3527_ (.A_N(_0546_),
    .B(_0557_),
    .C(_0558_),
    .D(\core_0.execute.rf.reg_outputs[3][5] ),
    .X(_0624_));
 sky130_fd_sc_hd__and4_1 _3528_ (.A(\core_0.execute.rf.reg_outputs[7][5] ),
    .B(_0546_),
    .C(_0530_),
    .D(_0531_),
    .X(_0625_));
 sky130_fd_sc_hd__a2111o_1 _3529_ (.A1(\core_0.execute.rf.reg_outputs[2][5] ),
    .A2(_0526_),
    .B1(_0624_),
    .C1(_0625_),
    .D1(_0566_),
    .X(_0626_));
 sky130_fd_sc_hd__o32ai_4 _3530_ (.A1(_0622_),
    .A2(_0623_),
    .A3(_0626_),
    .B1(_0521_),
    .B2(net99),
    .Y(_0627_));
 sky130_fd_sc_hd__clkinv_4 _3531_ (.A(_0627_),
    .Y(net205));
 sky130_fd_sc_hd__a22o_1 _3532_ (.A1(\core_0.execute.rf.reg_outputs[5][4] ),
    .A2(_0550_),
    .B1(_0555_),
    .B2(\core_0.execute.rf.reg_outputs[4][4] ),
    .X(_0628_));
 sky130_fd_sc_hd__a22o_1 _3533_ (.A1(\core_0.execute.rf.reg_outputs[1][4] ),
    .A2(_0542_),
    .B1(_0581_),
    .B2(\core_0.execute.rf.reg_outputs[6][4] ),
    .X(_0629_));
 sky130_fd_sc_hd__and4b_1 _3534_ (.A_N(_0546_),
    .B(_0530_),
    .C(_0531_),
    .D(\core_0.execute.rf.reg_outputs[3][4] ),
    .X(_0630_));
 sky130_fd_sc_hd__and4_1 _3535_ (.A(\core_0.execute.rf.reg_outputs[7][4] ),
    .B(_0546_),
    .C(_0530_),
    .D(_0531_),
    .X(_0631_));
 sky130_fd_sc_hd__a2111o_1 _3536_ (.A1(\core_0.execute.rf.reg_outputs[2][4] ),
    .A2(_0526_),
    .B1(_0630_),
    .C1(_0631_),
    .D1(_0566_),
    .X(_0632_));
 sky130_fd_sc_hd__o32ai_4 _3537_ (.A1(_0628_),
    .A2(_0629_),
    .A3(_0632_),
    .B1(_0521_),
    .B2(net98),
    .Y(_0633_));
 sky130_fd_sc_hd__clkinv_4 _3538_ (.A(_0633_),
    .Y(net204));
 sky130_fd_sc_hd__a22o_1 _3539_ (.A1(\core_0.execute.rf.reg_outputs[5][3] ),
    .A2(_0550_),
    .B1(_0555_),
    .B2(\core_0.execute.rf.reg_outputs[4][3] ),
    .X(_0634_));
 sky130_fd_sc_hd__a22o_1 _3540_ (.A1(\core_0.execute.rf.reg_outputs[3][3] ),
    .A2(_0522_),
    .B1(_0542_),
    .B2(\core_0.execute.rf.reg_outputs[1][3] ),
    .X(_0635_));
 sky130_fd_sc_hd__and4b_1 _3541_ (.A_N(_0518_),
    .B(_0537_),
    .C(_0523_),
    .D(\core_0.execute.rf.reg_outputs[6][3] ),
    .X(_0636_));
 sky130_fd_sc_hd__and4_1 _3542_ (.A(\core_0.execute.rf.reg_outputs[7][3] ),
    .B(_0523_),
    .C(_0517_),
    .D(_0524_),
    .X(_0637_));
 sky130_fd_sc_hd__a2111o_1 _3543_ (.A1(\core_0.execute.rf.reg_outputs[2][3] ),
    .A2(_0525_),
    .B1(_0636_),
    .C1(_0637_),
    .D1(_0566_),
    .X(_0638_));
 sky130_fd_sc_hd__o32ai_4 _3544_ (.A1(_0634_),
    .A2(_0635_),
    .A3(_0638_),
    .B1(_0520_),
    .B2(net97),
    .Y(_0639_));
 sky130_fd_sc_hd__inv_6 _3545_ (.A(_0639_),
    .Y(net203));
 sky130_fd_sc_hd__and2_1 _3546_ (.A(\core_0.execute.rf.reg_outputs[6][2] ),
    .B(_0581_),
    .X(_0640_));
 sky130_fd_sc_hd__a22o_1 _3547_ (.A1(\core_0.execute.rf.reg_outputs[7][2] ),
    .A2(_0545_),
    .B1(_0526_),
    .B2(\core_0.execute.rf.reg_outputs[2][2] ),
    .X(_0641_));
 sky130_fd_sc_hd__or2b_1 _3548_ (.A(\core_0.execute.rf.reg_outputs[4][2] ),
    .B_N(_0516_),
    .X(_0642_));
 sky130_fd_sc_hd__and4bb_1 _3549_ (.A_N(_0516_),
    .B_N(_0517_),
    .C(_0518_),
    .D(\core_0.execute.rf.reg_outputs[1][2] ),
    .X(_0643_));
 sky130_fd_sc_hd__and4b_1 _3550_ (.A_N(_0538_),
    .B(_0518_),
    .C(\core_0.execute.rf.reg_outputs[5][2] ),
    .D(_0516_),
    .X(_0644_));
 sky130_fd_sc_hd__and4b_1 _3551_ (.A_N(_0536_),
    .B(_0538_),
    .C(_0527_),
    .D(\core_0.execute.rf.reg_outputs[3][2] ),
    .X(_0645_));
 sky130_fd_sc_hd__a2111o_1 _3552_ (.A1(_0532_),
    .A2(_0642_),
    .B1(_0643_),
    .C1(_0644_),
    .D1(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__o32a_4 _3553_ (.A1(_0640_),
    .A2(_0641_),
    .A3(_0646_),
    .B1(_0520_),
    .B2(net96),
    .X(_0647_));
 sky130_fd_sc_hd__buf_8 _3554_ (.A(_0647_),
    .X(net202));
 sky130_fd_sc_hd__and4b_1 _3555_ (.A_N(_0557_),
    .B(_0527_),
    .C(\core_0.execute.rf.reg_outputs[5][1] ),
    .D(_0536_),
    .X(_0648_));
 sky130_fd_sc_hd__and4bb_1 _3556_ (.A_N(_0556_),
    .B_N(_0557_),
    .C(_0558_),
    .D(\core_0.execute.rf.reg_outputs[1][1] ),
    .X(_0649_));
 sky130_fd_sc_hd__and4b_1 _3557_ (.A_N(_0546_),
    .B(_0557_),
    .C(_0558_),
    .D(\core_0.execute.rf.reg_outputs[3][1] ),
    .X(_0650_));
 sky130_fd_sc_hd__a2111o_4 _3558_ (.A1(\core_0.execute.rf.reg_outputs[4][1] ),
    .A2(_0555_),
    .B1(_0648_),
    .C1(_0649_),
    .D1(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__and4_1 _3559_ (.A(\core_0.execute.rf.reg_outputs[7][1] ),
    .B(_0536_),
    .C(_0538_),
    .D(_0527_),
    .X(_0652_));
 sky130_fd_sc_hd__and4b_1 _3560_ (.A_N(_0558_),
    .B(_0538_),
    .C(_0556_),
    .D(\core_0.execute.rf.reg_outputs[6][1] ),
    .X(_0653_));
 sky130_fd_sc_hd__a2111o_4 _3561_ (.A1(\core_0.execute.rf.reg_outputs[2][1] ),
    .A2(_0526_),
    .B1(_0652_),
    .C1(_0653_),
    .D1(_0566_),
    .X(_0654_));
 sky130_fd_sc_hd__o22ai_4 _3562_ (.A1(net95),
    .A2(_0521_),
    .B1(_0651_),
    .B2(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__clkinv_4 _3563_ (.A(_0655_),
    .Y(net201));
 sky130_fd_sc_hd__and4b_1 _3564_ (.A_N(_0571_),
    .B(_0569_),
    .C(_0573_),
    .D(\core_0.execute.rf.reg_outputs[6][0] ),
    .X(_0656_));
 sky130_fd_sc_hd__and4bb_1 _3565_ (.A_N(_0573_),
    .B_N(_0571_),
    .C(_0569_),
    .D(\core_0.execute.rf.reg_outputs[2][0] ),
    .X(_0657_));
 sky130_fd_sc_hd__and4b_1 _3566_ (.A_N(_0573_),
    .B(_0569_),
    .C(_0571_),
    .D(\core_0.execute.rf.reg_outputs[3][0] ),
    .X(_0658_));
 sky130_fd_sc_hd__a2111oi_4 _3567_ (.A1(\core_0.execute.rf.reg_outputs[1][0] ),
    .A2(_0542_),
    .B1(_0656_),
    .C1(_0657_),
    .D1(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__and4_1 _3568_ (.A(\core_0.execute.rf.reg_outputs[7][0] ),
    .B(_0573_),
    .C(_0569_),
    .D(_0571_),
    .X(_0660_));
 sky130_fd_sc_hd__and4b_1 _3569_ (.A_N(_0569_),
    .B(_0571_),
    .C(\core_0.execute.rf.reg_outputs[5][0] ),
    .D(_0573_),
    .X(_0661_));
 sky130_fd_sc_hd__a2111oi_4 _3570_ (.A1(\core_0.execute.rf.reg_outputs[4][0] ),
    .A2(_0555_),
    .B1(_0660_),
    .C1(_0661_),
    .D1(_0566_),
    .Y(_0662_));
 sky130_fd_sc_hd__nor2_2 _3571_ (.A(net88),
    .B(_0521_),
    .Y(_0663_));
 sky130_fd_sc_hd__a21o_4 _3572_ (.A1(_0659_),
    .A2(_0662_),
    .B1(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__clkinv_4 _3573_ (.A(_0664_),
    .Y(net194));
 sky130_fd_sc_hd__clkinv_2 _3574_ (.A(net71),
    .Y(_0665_));
 sky130_fd_sc_hd__inv_2 _3575_ (.A(\core_0.fetch.dbg_out ),
    .Y(_0666_));
 sky130_fd_sc_hd__clkbuf_4 _3576_ (.A(\core_0.fetch.out_buffer_valid ),
    .X(_0667_));
 sky130_fd_sc_hd__buf_6 _3577_ (.A(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__buf_4 _3578_ (.A(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__buf_4 _3579_ (.A(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__o21a_1 _3580_ (.A1(net19),
    .A2(net18),
    .B1(\core_0.execute.irq_en ),
    .X(_0671_));
 sky130_fd_sc_hd__or3_1 _3581_ (.A(net37),
    .B(\core_0.execute.sreg_irq_flags.i_d[2] ),
    .C(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__or2_1 _3582_ (.A(\core_0.execute.prev_sys ),
    .B(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__buf_4 _3583_ (.A(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__buf_6 _3584_ (.A(net105),
    .X(_0675_));
 sky130_fd_sc_hd__nand2_4 _3585_ (.A(\core_0.execute.pc_high_out[2] ),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__nand2_4 _3586_ (.A(\core_0.execute.pc_high_out[7] ),
    .B(_0675_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand2_4 _3587_ (.A(\core_0.execute.pc_high_out[3] ),
    .B(_0675_),
    .Y(_0678_));
 sky130_fd_sc_hd__a2bb2o_1 _3588_ (.A1_N(\core_0.execute.prev_pc_high[7] ),
    .A2_N(_0677_),
    .B1(_0678_),
    .B2(\core_0.execute.prev_pc_high[3] ),
    .X(_0679_));
 sky130_fd_sc_hd__a221o_1 _3589_ (.A1(\core_0.execute.prev_pc_high[2] ),
    .A2(_0676_),
    .B1(_0677_),
    .B2(\core_0.execute.prev_pc_high[7] ),
    .C1(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__nand2_4 _3590_ (.A(\core_0.execute.pc_high_out[6] ),
    .B(_0675_),
    .Y(_0681_));
 sky130_fd_sc_hd__nand2_4 _3591_ (.A(\core_0.execute.pc_high_out[4] ),
    .B(net105),
    .Y(_0682_));
 sky130_fd_sc_hd__o2bb2a_1 _3592_ (.A1_N(\core_0.execute.prev_pc_high[6] ),
    .A2_N(_0681_),
    .B1(_0682_),
    .B2(\core_0.execute.prev_pc_high[4] ),
    .X(_0683_));
 sky130_fd_sc_hd__o221ai_1 _3593_ (.A1(\core_0.execute.prev_pc_high[6] ),
    .A2(_0681_),
    .B1(_0676_),
    .B2(\core_0.execute.prev_pc_high[2] ),
    .C1(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2_4 _3594_ (.A(\core_0.execute.pc_high_out[5] ),
    .B(net105),
    .Y(_0685_));
 sky130_fd_sc_hd__xnor2_1 _3595_ (.A(\core_0.execute.prev_pc_high[5] ),
    .B(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__nand2_2 _3596_ (.A(\core_0.execute.pc_high_out[1] ),
    .B(net105),
    .Y(_0687_));
 sky130_fd_sc_hd__a2bb2o_1 _3597_ (.A1_N(\core_0.execute.prev_pc_high[1] ),
    .A2_N(_0687_),
    .B1(_0682_),
    .B2(\core_0.execute.prev_pc_high[4] ),
    .X(_0688_));
 sky130_fd_sc_hd__nand2_2 _3598_ (.A(\core_0.execute.pc_high_out[0] ),
    .B(_0675_),
    .Y(_0689_));
 sky130_fd_sc_hd__xnor2_1 _3599_ (.A(\core_0.execute.prev_pc_high[0] ),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__a2bb2o_1 _3600_ (.A1_N(\core_0.execute.prev_pc_high[3] ),
    .A2_N(_0678_),
    .B1(_0687_),
    .B2(\core_0.execute.prev_pc_high[1] ),
    .X(_0691_));
 sky130_fd_sc_hd__or4_1 _3601_ (.A(_0686_),
    .B(_0688_),
    .C(_0690_),
    .D(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__or3_2 _3602_ (.A(_0680_),
    .B(_0684_),
    .C(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__or2_2 _3603_ (.A(_0674_),
    .B(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__nor2_1 _3604_ (.A(\core_0.execute.hold_valid ),
    .B(\core_0.decode.o_submit ),
    .Y(_0695_));
 sky130_fd_sc_hd__or3_1 _3605_ (.A(\core_0.decode.i_flush ),
    .B(_0694_),
    .C(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__clkbuf_4 _3606_ (.A(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__inv_2 _3607_ (.A(\core_0.execute.next_ready_delayed ),
    .Y(_0698_));
 sky130_fd_sc_hd__clkbuf_4 _3608_ (.A(\core_0.dec_l_reg_sel[2] ),
    .X(_0699_));
 sky130_fd_sc_hd__buf_2 _3609_ (.A(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__buf_2 _3610_ (.A(\core_0.dec_l_reg_sel[1] ),
    .X(_0701_));
 sky130_fd_sc_hd__clkbuf_4 _3611_ (.A(\core_0.dec_l_reg_sel[0] ),
    .X(_0702_));
 sky130_fd_sc_hd__and3_4 _3612_ (.A(_0700_),
    .B(_0701_),
    .C(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__clkbuf_4 _3613_ (.A(_0701_),
    .X(_0704_));
 sky130_fd_sc_hd__inv_2 _3614_ (.A(_0702_),
    .Y(_0705_));
 sky130_fd_sc_hd__clkbuf_4 _3615_ (.A(_0700_),
    .X(_0706_));
 sky130_fd_sc_hd__a31o_1 _3616_ (.A1(_0704_),
    .A2(_0705_),
    .A3(\core_0.ew_reg_ie[3] ),
    .B1(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__buf_4 _3617_ (.A(\core_0.dec_l_reg_sel[1] ),
    .X(_0708_));
 sky130_fd_sc_hd__clkbuf_4 _3618_ (.A(\core_0.dec_l_reg_sel[0] ),
    .X(_0709_));
 sky130_fd_sc_hd__nor2_2 _3619_ (.A(_0708_),
    .B(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__buf_4 _3620_ (.A(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__or2_1 _3621_ (.A(_0704_),
    .B(\core_0.ew_reg_ie[2] ),
    .X(_0712_));
 sky130_fd_sc_hd__clkbuf_4 _3622_ (.A(_0702_),
    .X(_0713_));
 sky130_fd_sc_hd__buf_4 _3623_ (.A(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__buf_4 _3624_ (.A(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__a22o_1 _3625_ (.A1(\core_0.ew_reg_ie[1] ),
    .A2(_0711_),
    .B1(_0712_),
    .B2(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__inv_2 _3626_ (.A(_0700_),
    .Y(_0717_));
 sky130_fd_sc_hd__nand2_1 _3627_ (.A(_0704_),
    .B(_0715_),
    .Y(_0718_));
 sky130_fd_sc_hd__and2_1 _3628_ (.A(_0717_),
    .B(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__mux4_1 _3629_ (.A0(\core_0.ew_reg_ie[5] ),
    .A1(\core_0.ew_reg_ie[6] ),
    .A2(\core_0.ew_reg_ie[7] ),
    .A3(\core_0.ew_reg_ie[4] ),
    .S0(_0715_),
    .S1(_0704_),
    .X(_0720_));
 sky130_fd_sc_hd__and2_1 _3630_ (.A(\core_0.execute.sreg_long_ptr_en ),
    .B(\core_0.dec_mem_long ),
    .X(_0721_));
 sky130_fd_sc_hd__o21a_1 _3631_ (.A1(_0719_),
    .A2(_0720_),
    .B1(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__o21ai_1 _3632_ (.A1(_0707_),
    .A2(_0716_),
    .B1(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__mux2_1 _3633_ (.A0(\core_0.ew_reg_ie[0] ),
    .A1(\core_0.ew_reg_ie[1] ),
    .S(_0715_),
    .X(_0724_));
 sky130_fd_sc_hd__nand2_1 _3634_ (.A(_0704_),
    .B(_0705_),
    .Y(_0725_));
 sky130_fd_sc_hd__o221a_1 _3635_ (.A1(\core_0.ew_reg_ie[2] ),
    .A2(_0725_),
    .B1(_0718_),
    .B2(\core_0.ew_reg_ie[3] ),
    .C1(_0717_),
    .X(_0726_));
 sky130_fd_sc_hd__o21ai_1 _3636_ (.A1(_0704_),
    .A2(_0724_),
    .B1(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__mux2_1 _3637_ (.A0(\core_0.ew_reg_ie[4] ),
    .A1(\core_0.ew_reg_ie[5] ),
    .S(_0715_),
    .X(_0728_));
 sky130_fd_sc_hd__o221a_1 _3638_ (.A1(\core_0.ew_reg_ie[6] ),
    .A2(_0725_),
    .B1(_0718_),
    .B2(\core_0.ew_reg_ie[7] ),
    .C1(_0706_),
    .X(_0729_));
 sky130_fd_sc_hd__o21ai_1 _3639_ (.A1(_0704_),
    .A2(_0728_),
    .B1(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__o211a_1 _3640_ (.A1(_0703_),
    .A2(_0723_),
    .B1(_0727_),
    .C1(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__and2b_1 _3641_ (.A_N(_0731_),
    .B(\core_0.dec_used_operands[0] ),
    .X(_0732_));
 sky130_fd_sc_hd__mux4_1 _3642_ (.A0(\core_0.ew_reg_ie[0] ),
    .A1(\core_0.ew_reg_ie[1] ),
    .A2(\core_0.ew_reg_ie[2] ),
    .A3(\core_0.ew_reg_ie[3] ),
    .S0(_0571_),
    .S1(_0569_),
    .X(_0733_));
 sky130_fd_sc_hd__clkinv_2 _3643_ (.A(_0573_),
    .Y(_0734_));
 sky130_fd_sc_hd__mux4_1 _3644_ (.A0(\core_0.ew_reg_ie[4] ),
    .A1(\core_0.ew_reg_ie[5] ),
    .A2(\core_0.ew_reg_ie[6] ),
    .A3(\core_0.ew_reg_ie[7] ),
    .S0(_0571_),
    .S1(_0569_),
    .X(_0735_));
 sky130_fd_sc_hd__or2_1 _3645_ (.A(_0734_),
    .B(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__o211a_1 _3646_ (.A1(_0573_),
    .A2(_0733_),
    .B1(_0736_),
    .C1(\core_0.dec_used_operands[1] ),
    .X(_0737_));
 sky130_fd_sc_hd__o22a_2 _3647_ (.A1(\core_0.ew_submit ),
    .A2(_0698_),
    .B1(_0732_),
    .B2(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__inv_2 _3648_ (.A(net20),
    .Y(_0739_));
 sky130_fd_sc_hd__a22o_4 _3649_ (.A1(net156),
    .A2(_0739_),
    .B1(\core_0.ew_mem_access ),
    .B2(\core_0.ew_submit ),
    .X(_0740_));
 sky130_fd_sc_hd__or2_4 _3650_ (.A(\core_0.execute.alu_mul_div.i_div ),
    .B(\core_0.execute.alu_mul_div.i_mod ),
    .X(_0741_));
 sky130_fd_sc_hd__nand2_4 _3651_ (.A(\core_0.decode.o_submit ),
    .B(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__nand2_4 _3652_ (.A(\core_0.decode.o_submit ),
    .B(\core_0.execute.alu_mul_div.i_mul ),
    .Y(_0743_));
 sky130_fd_sc_hd__nand2_2 _3653_ (.A(_0742_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__or3_2 _3654_ (.A(\core_0.execute.alu_mul_div.comp ),
    .B(_0740_),
    .C(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__nor3_4 _3655_ (.A(_0738_),
    .B(_0745_),
    .C(_0696_),
    .Y(_0746_));
 sky130_fd_sc_hd__nor2_4 _3656_ (.A(_0697_),
    .B(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__nor2_4 _3657_ (.A(\core_0.decode.input_valid ),
    .B(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__mux2_1 _3658_ (.A0(net66),
    .A1(\core_0.fetch.out_buffer_data_instr[6] ),
    .S(_0669_),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _3659_ (.A0(net65),
    .A1(\core_0.fetch.out_buffer_data_instr[5] ),
    .S(_0669_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_2 _3660_ (.A0(net38),
    .A1(\core_0.fetch.out_buffer_data_instr[0] ),
    .S(_0668_),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_2 _3661_ (.A0(net49),
    .A1(\core_0.fetch.out_buffer_data_instr[1] ),
    .S(_0668_),
    .X(_0752_));
 sky130_fd_sc_hd__or2b_1 _3662_ (.A(_0751_),
    .B_N(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _3663_ (.A0(net60),
    .A1(\core_0.fetch.out_buffer_data_instr[2] ),
    .S(_0669_),
    .X(_0754_));
 sky130_fd_sc_hd__mux2_1 _3664_ (.A0(net63),
    .A1(\core_0.fetch.out_buffer_data_instr[3] ),
    .S(_0669_),
    .X(_0755_));
 sky130_fd_sc_hd__nand2_1 _3665_ (.A(_0754_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__nor2_1 _3666_ (.A(_0753_),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__mux2_2 _3667_ (.A0(net54),
    .A1(\core_0.fetch.out_buffer_data_instr[24] ),
    .S(_0668_),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_2 _3668_ (.A0(net46),
    .A1(\core_0.fetch.out_buffer_data_instr[17] ),
    .S(\core_0.fetch.out_buffer_valid ),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_4 _3669_ (.A0(net56),
    .A1(\core_0.fetch.out_buffer_data_instr[26] ),
    .S(_0668_),
    .X(_0760_));
 sky130_fd_sc_hd__mux2_2 _3670_ (.A0(net48),
    .A1(\core_0.fetch.out_buffer_data_instr[19] ),
    .S(\core_0.fetch.out_buffer_valid ),
    .X(_0761_));
 sky130_fd_sc_hd__or4_1 _3671_ (.A(_0758_),
    .B(_0759_),
    .C(_0760_),
    .D(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__mux2_2 _3672_ (.A0(net50),
    .A1(\core_0.fetch.out_buffer_data_instr[20] ),
    .S(\core_0.fetch.out_buffer_valid ),
    .X(_0763_));
 sky130_fd_sc_hd__mux2_2 _3673_ (.A0(net61),
    .A1(\core_0.fetch.out_buffer_data_instr[30] ),
    .S(_0667_),
    .X(_0764_));
 sky130_fd_sc_hd__mux2_4 _3674_ (.A0(net53),
    .A1(\core_0.fetch.out_buffer_data_instr[23] ),
    .S(_0667_),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_2 _3675_ (.A0(net47),
    .A1(\core_0.fetch.out_buffer_data_instr[18] ),
    .S(\core_0.fetch.out_buffer_valid ),
    .X(_0766_));
 sky130_fd_sc_hd__or4_1 _3676_ (.A(_0763_),
    .B(_0764_),
    .C(_0765_),
    .D(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_2 _3677_ (.A0(net58),
    .A1(\core_0.fetch.out_buffer_data_instr[28] ),
    .S(_0667_),
    .X(_0768_));
 sky130_fd_sc_hd__or2b_1 _3678_ (.A(\core_0.fetch.out_buffer_data_instr[31] ),
    .B_N(_0667_),
    .X(_0769_));
 sky130_fd_sc_hd__o21a_1 _3679_ (.A1(_0668_),
    .A2(net62),
    .B1(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__mux2_2 _3680_ (.A0(net45),
    .A1(\core_0.fetch.out_buffer_data_instr[16] ),
    .S(\core_0.fetch.out_buffer_valid ),
    .X(_0771_));
 sky130_fd_sc_hd__mux2_2 _3681_ (.A0(net51),
    .A1(\core_0.fetch.out_buffer_data_instr[21] ),
    .S(_0667_),
    .X(_0772_));
 sky130_fd_sc_hd__or4_1 _3682_ (.A(_0768_),
    .B(_0770_),
    .C(_0771_),
    .D(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_2 _3683_ (.A0(net52),
    .A1(\core_0.fetch.out_buffer_data_instr[22] ),
    .S(_0667_),
    .X(_0774_));
 sky130_fd_sc_hd__or2b_1 _3684_ (.A(\core_0.fetch.out_buffer_data_instr[27] ),
    .B_N(_0667_),
    .X(_0775_));
 sky130_fd_sc_hd__o21a_1 _3685_ (.A1(_0668_),
    .A2(net57),
    .B1(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__or2b_1 _3686_ (.A(\core_0.fetch.out_buffer_data_instr[25] ),
    .B_N(_0667_),
    .X(_0777_));
 sky130_fd_sc_hd__o21a_1 _3687_ (.A1(_0668_),
    .A2(net55),
    .B1(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_2 _3688_ (.A0(net59),
    .A1(\core_0.fetch.out_buffer_data_instr[29] ),
    .S(_0667_),
    .X(_0779_));
 sky130_fd_sc_hd__or4_1 _3689_ (.A(_0774_),
    .B(_0776_),
    .C(_0778_),
    .D(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__or3_2 _3690_ (.A(_0767_),
    .B(_0773_),
    .C(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__or4b_1 _3691_ (.A(_0752_),
    .B(_0762_),
    .C(_0781_),
    .D_N(_0751_),
    .X(_0782_));
 sky130_fd_sc_hd__a211oi_1 _3692_ (.A1(_0753_),
    .A2(_0782_),
    .B1(_0754_),
    .C1(_0755_),
    .Y(_0783_));
 sky130_fd_sc_hd__nor2_1 _3693_ (.A(_0757_),
    .B(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__mux2_1 _3694_ (.A0(net64),
    .A1(\core_0.fetch.out_buffer_data_instr[4] ),
    .S(_0669_),
    .X(_0785_));
 sky130_fd_sc_hd__or4b_1 _3695_ (.A(_0749_),
    .B(_0750_),
    .C(_0784_),
    .D_N(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__o211a_1 _3696_ (.A1(_0670_),
    .A2(net70),
    .B1(_0748_),
    .C1(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__a211o_4 _3697_ (.A1(\core_0.fetch.pc_flush_override ),
    .A2(_0666_),
    .B1(_0787_),
    .C1(\core_0.fetch.pc_reset_override ),
    .X(_0788_));
 sky130_fd_sc_hd__and2_1 _3698_ (.A(_0665_),
    .B(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__clkbuf_4 _3699_ (.A(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__buf_6 _3700_ (.A(_0790_),
    .X(net177));
 sky130_fd_sc_hd__buf_6 _3701_ (.A(\core_0.decode.i_flush ),
    .X(_0791_));
 sky130_fd_sc_hd__nor2_2 _3702_ (.A(\core_0.fetch.pc_flush_override ),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__clkbuf_4 _3703_ (.A(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__inv_2 _3704_ (.A(\core_0.fetch.prev_request_pc[14] ),
    .Y(_0794_));
 sky130_fd_sc_hd__o21ai_1 _3705_ (.A1(_0669_),
    .A2(net62),
    .B1(_0769_),
    .Y(_0795_));
 sky130_fd_sc_hd__o2bb2a_1 _3706_ (.A1_N(_0764_),
    .A2_N(_0794_),
    .B1(\core_0.fetch.prev_request_pc[15] ),
    .B2(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__inv_2 _3707_ (.A(\core_0.fetch.prev_request_pc[12] ),
    .Y(_0797_));
 sky130_fd_sc_hd__inv_2 _3708_ (.A(\core_0.fetch.prev_request_pc[13] ),
    .Y(_0798_));
 sky130_fd_sc_hd__o21ai_2 _3709_ (.A1(_0668_),
    .A2(net57),
    .B1(_0775_),
    .Y(_0799_));
 sky130_fd_sc_hd__inv_2 _3710_ (.A(\core_0.fetch.prev_request_pc[10] ),
    .Y(_0800_));
 sky130_fd_sc_hd__a2bb2o_1 _3711_ (.A1_N(\core_0.fetch.prev_request_pc[11] ),
    .A2_N(_0799_),
    .B1(_0760_),
    .B2(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__nand2_1 _3712_ (.A(\core_0.fetch.prev_request_pc[11] ),
    .B(_0799_),
    .Y(_0802_));
 sky130_fd_sc_hd__o21ai_1 _3713_ (.A1(_0800_),
    .A2(_0760_),
    .B1(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__nor2_1 _3714_ (.A(_0801_),
    .B(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__inv_2 _3715_ (.A(\core_0.fetch.prev_request_pc[6] ),
    .Y(_0805_));
 sky130_fd_sc_hd__inv_2 _3716_ (.A(\core_0.fetch.prev_request_pc[7] ),
    .Y(_0806_));
 sky130_fd_sc_hd__inv_2 _3717_ (.A(\core_0.fetch.prev_request_pc[5] ),
    .Y(_0807_));
 sky130_fd_sc_hd__inv_2 _3718_ (.A(\core_0.fetch.prev_request_pc[4] ),
    .Y(_0808_));
 sky130_fd_sc_hd__inv_2 _3719_ (.A(\core_0.fetch.prev_request_pc[3] ),
    .Y(_0809_));
 sky130_fd_sc_hd__inv_2 _3720_ (.A(\core_0.fetch.prev_request_pc[2] ),
    .Y(_0810_));
 sky130_fd_sc_hd__inv_2 _3721_ (.A(\core_0.fetch.prev_request_pc[1] ),
    .Y(_0811_));
 sky130_fd_sc_hd__inv_2 _3722_ (.A(\core_0.fetch.prev_request_pc[0] ),
    .Y(_0812_));
 sky130_fd_sc_hd__a211o_1 _3723_ (.A1(_0811_),
    .A2(_0759_),
    .B1(_0771_),
    .C1(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__o221a_1 _3724_ (.A1(_0811_),
    .A2(_0759_),
    .B1(_0766_),
    .B2(_0810_),
    .C1(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__a221o_1 _3725_ (.A1(_0809_),
    .A2(_0761_),
    .B1(_0766_),
    .B2(_0810_),
    .C1(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__o221a_1 _3726_ (.A1(_0808_),
    .A2(_0763_),
    .B1(_0761_),
    .B2(_0809_),
    .C1(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__a221o_1 _3727_ (.A1(_0808_),
    .A2(_0763_),
    .B1(_0772_),
    .B2(_0807_),
    .C1(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__o221a_1 _3728_ (.A1(_0805_),
    .A2(_0774_),
    .B1(_0772_),
    .B2(_0807_),
    .C1(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__a221o_1 _3729_ (.A1(_0805_),
    .A2(_0774_),
    .B1(_0765_),
    .B2(_0806_),
    .C1(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__o21ai_2 _3730_ (.A1(_0668_),
    .A2(net55),
    .B1(_0777_),
    .Y(_0820_));
 sky130_fd_sc_hd__inv_2 _3731_ (.A(\core_0.fetch.prev_request_pc[8] ),
    .Y(_0821_));
 sky130_fd_sc_hd__a2bb2o_1 _3732_ (.A1_N(\core_0.fetch.prev_request_pc[9] ),
    .A2_N(_0820_),
    .B1(_0758_),
    .B2(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__nand2_1 _3733_ (.A(\core_0.fetch.prev_request_pc[9] ),
    .B(_0820_),
    .Y(_0823_));
 sky130_fd_sc_hd__o221a_1 _3734_ (.A1(_0821_),
    .A2(_0758_),
    .B1(_0765_),
    .B2(_0806_),
    .C1(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__and2b_1 _3735_ (.A_N(_0822_),
    .B(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__a32o_1 _3736_ (.A1(_0804_),
    .A2(_0823_),
    .A3(_0822_),
    .B1(_0802_),
    .B2(_0801_),
    .X(_0826_));
 sky130_fd_sc_hd__a31o_1 _3737_ (.A1(_0804_),
    .A2(_0819_),
    .A3(_0825_),
    .B1(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__o21a_1 _3738_ (.A1(_0797_),
    .A2(_0768_),
    .B1(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__a221o_1 _3739_ (.A1(_0797_),
    .A2(_0768_),
    .B1(_0779_),
    .B2(_0798_),
    .C1(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__nand2_1 _3740_ (.A(\core_0.fetch.prev_request_pc[15] ),
    .B(_0795_),
    .Y(_0830_));
 sky130_fd_sc_hd__o221a_1 _3741_ (.A1(_0794_),
    .A2(_0764_),
    .B1(_0779_),
    .B2(_0798_),
    .C1(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__and2b_1 _3742_ (.A_N(_0796_),
    .B(_0830_),
    .X(_0832_));
 sky130_fd_sc_hd__a31o_1 _3743_ (.A1(_0796_),
    .A2(_0829_),
    .A3(_0831_),
    .B1(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_1 _3744_ (.A0(net69),
    .A1(\core_0.fetch.out_buffer_data_instr[9] ),
    .S(_0669_),
    .X(_0834_));
 sky130_fd_sc_hd__mux2_1 _3745_ (.A0(net67),
    .A1(\core_0.fetch.out_buffer_data_instr[7] ),
    .S(_0669_),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _3746_ (.A0(net39),
    .A1(\core_0.fetch.out_buffer_data_instr[10] ),
    .S(_0669_),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_1 _3747_ (.A0(net68),
    .A1(\core_0.fetch.out_buffer_data_instr[8] ),
    .S(_0670_),
    .X(_0837_));
 sky130_fd_sc_hd__o41a_1 _3748_ (.A1(_0834_),
    .A2(_0835_),
    .A3(_0836_),
    .A4(_0837_),
    .B1(_0757_),
    .X(_0838_));
 sky130_fd_sc_hd__or3_1 _3749_ (.A(_0749_),
    .B(_0750_),
    .C(_0756_),
    .X(_0839_));
 sky130_fd_sc_hd__or4b_1 _3750_ (.A(\core_0.fetch.pc_reset_override ),
    .B(_0785_),
    .C(_0839_),
    .D_N(_0752_),
    .X(_0840_));
 sky130_fd_sc_hd__a21oi_1 _3751_ (.A1(_0833_),
    .A2(_0838_),
    .B1(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__clkbuf_4 _3752_ (.A(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__or2_4 _3753_ (.A(\core_0.fetch.pc_flush_override ),
    .B(_0791_),
    .X(_0843_));
 sky130_fd_sc_hd__a21o_1 _3754_ (.A1(_0770_),
    .A2(_0842_),
    .B1(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__clkbuf_4 _3755_ (.A(_0842_),
    .X(_0845_));
 sky130_fd_sc_hd__and3_1 _3756_ (.A(\core_0.fetch.prev_request_pc[2] ),
    .B(\core_0.fetch.prev_request_pc[1] ),
    .C(\core_0.fetch.prev_request_pc[0] ),
    .X(_0846_));
 sky130_fd_sc_hd__and2_1 _3757_ (.A(\core_0.fetch.prev_request_pc[3] ),
    .B(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__and3_1 _3758_ (.A(\core_0.fetch.prev_request_pc[5] ),
    .B(\core_0.fetch.prev_request_pc[4] ),
    .C(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__and3_1 _3759_ (.A(\core_0.fetch.prev_request_pc[7] ),
    .B(\core_0.fetch.prev_request_pc[6] ),
    .C(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__and2_1 _3760_ (.A(\core_0.fetch.prev_request_pc[8] ),
    .B(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__and3_1 _3761_ (.A(\core_0.fetch.prev_request_pc[10] ),
    .B(\core_0.fetch.prev_request_pc[9] ),
    .C(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__and2_1 _3762_ (.A(\core_0.fetch.prev_request_pc[11] ),
    .B(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__and3_1 _3763_ (.A(\core_0.fetch.prev_request_pc[13] ),
    .B(\core_0.fetch.prev_request_pc[12] ),
    .C(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__and2_1 _3764_ (.A(\core_0.fetch.prev_request_pc[14] ),
    .B(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__xnor2_1 _3765_ (.A(\core_0.fetch.prev_request_pc[15] ),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__nor2_1 _3766_ (.A(_0845_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__clkinv_2 _3767_ (.A(\core_0.fetch.pc_reset_override ),
    .Y(_0857_));
 sky130_fd_sc_hd__clkbuf_4 _3768_ (.A(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__o221a_1 _3769_ (.A1(net78),
    .A2(_0793_),
    .B1(_0844_),
    .B2(_0856_),
    .C1(_0858_),
    .X(net167));
 sky130_fd_sc_hd__nor2_1 _3770_ (.A(\core_0.fetch.prev_request_pc[14] ),
    .B(_0853_),
    .Y(_0859_));
 sky130_fd_sc_hd__nor3_1 _3771_ (.A(_0845_),
    .B(_0854_),
    .C(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__clkbuf_4 _3772_ (.A(_0841_),
    .X(_0861_));
 sky130_fd_sc_hd__clkbuf_4 _3773_ (.A(_0843_),
    .X(_0862_));
 sky130_fd_sc_hd__a21o_1 _3774_ (.A1(_0764_),
    .A2(_0861_),
    .B1(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__o221a_1 _3775_ (.A1(net77),
    .A2(_0793_),
    .B1(_0860_),
    .B2(_0863_),
    .C1(_0858_),
    .X(net166));
 sky130_fd_sc_hd__a21oi_1 _3776_ (.A1(\core_0.fetch.prev_request_pc[12] ),
    .A2(_0852_),
    .B1(\core_0.fetch.prev_request_pc[13] ),
    .Y(_0864_));
 sky130_fd_sc_hd__nor3_1 _3777_ (.A(_0845_),
    .B(_0853_),
    .C(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__a21o_1 _3778_ (.A1(_0779_),
    .A2(_0861_),
    .B1(_0862_),
    .X(_0866_));
 sky130_fd_sc_hd__o221a_1 _3779_ (.A1(net76),
    .A2(_0793_),
    .B1(_0865_),
    .B2(_0866_),
    .C1(_0858_),
    .X(net165));
 sky130_fd_sc_hd__xnor2_1 _3780_ (.A(_0797_),
    .B(_0852_),
    .Y(_0867_));
 sky130_fd_sc_hd__mux2_1 _3781_ (.A0(_0867_),
    .A1(_0768_),
    .S(_0842_),
    .X(_0868_));
 sky130_fd_sc_hd__or2_1 _3782_ (.A(net75),
    .B(_0792_),
    .X(_0869_));
 sky130_fd_sc_hd__o211a_1 _3783_ (.A1(_0862_),
    .A2(_0868_),
    .B1(_0869_),
    .C1(_0858_),
    .X(net164));
 sky130_fd_sc_hd__nor2_1 _3784_ (.A(\core_0.fetch.prev_request_pc[11] ),
    .B(_0851_),
    .Y(_0870_));
 sky130_fd_sc_hd__nor3_1 _3785_ (.A(_0845_),
    .B(_0852_),
    .C(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__a21o_1 _3786_ (.A1(_0776_),
    .A2(_0861_),
    .B1(_0862_),
    .X(_0872_));
 sky130_fd_sc_hd__o221a_1 _3787_ (.A1(net74),
    .A2(_0793_),
    .B1(_0871_),
    .B2(_0872_),
    .C1(_0858_),
    .X(net163));
 sky130_fd_sc_hd__a21oi_1 _3788_ (.A1(\core_0.fetch.prev_request_pc[9] ),
    .A2(_0850_),
    .B1(\core_0.fetch.prev_request_pc[10] ),
    .Y(_0873_));
 sky130_fd_sc_hd__nor3_1 _3789_ (.A(_0845_),
    .B(_0851_),
    .C(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__a21o_1 _3790_ (.A1(_0760_),
    .A2(_0861_),
    .B1(_0862_),
    .X(_0875_));
 sky130_fd_sc_hd__o221a_1 _3791_ (.A1(net73),
    .A2(_0793_),
    .B1(_0874_),
    .B2(_0875_),
    .C1(_0858_),
    .X(net162));
 sky130_fd_sc_hd__xnor2_1 _3792_ (.A(\core_0.fetch.prev_request_pc[9] ),
    .B(_0850_),
    .Y(_0876_));
 sky130_fd_sc_hd__nor2_1 _3793_ (.A(_0842_),
    .B(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__a211o_1 _3794_ (.A1(_0778_),
    .A2(_0842_),
    .B1(_0843_),
    .C1(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__o211a_2 _3795_ (.A1(net87),
    .A2(_0793_),
    .B1(_0878_),
    .C1(_0858_),
    .X(net176));
 sky130_fd_sc_hd__nor2_1 _3796_ (.A(\core_0.fetch.prev_request_pc[8] ),
    .B(_0849_),
    .Y(_0879_));
 sky130_fd_sc_hd__nor2_1 _3797_ (.A(_0850_),
    .B(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__mux2_1 _3798_ (.A0(_0880_),
    .A1(_0758_),
    .S(_0842_),
    .X(_0881_));
 sky130_fd_sc_hd__or2_1 _3799_ (.A(net86),
    .B(_0792_),
    .X(_0882_));
 sky130_fd_sc_hd__o211a_1 _3800_ (.A1(_0862_),
    .A2(_0881_),
    .B1(_0882_),
    .C1(_0858_),
    .X(net175));
 sky130_fd_sc_hd__and2_1 _3801_ (.A(\core_0.fetch.prev_request_pc[6] ),
    .B(_0848_),
    .X(_0883_));
 sky130_fd_sc_hd__nor2_1 _3802_ (.A(\core_0.fetch.prev_request_pc[7] ),
    .B(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__nor3_1 _3803_ (.A(_0845_),
    .B(_0849_),
    .C(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__a21o_1 _3804_ (.A1(_0765_),
    .A2(_0861_),
    .B1(_0862_),
    .X(_0886_));
 sky130_fd_sc_hd__o221a_2 _3805_ (.A1(net85),
    .A2(_0793_),
    .B1(_0885_),
    .B2(_0886_),
    .C1(_0858_),
    .X(net174));
 sky130_fd_sc_hd__nor2_1 _3806_ (.A(\core_0.fetch.prev_request_pc[6] ),
    .B(_0848_),
    .Y(_0887_));
 sky130_fd_sc_hd__nor3_1 _3807_ (.A(_0845_),
    .B(_0883_),
    .C(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__a21o_1 _3808_ (.A1(_0774_),
    .A2(_0861_),
    .B1(_0862_),
    .X(_0889_));
 sky130_fd_sc_hd__o221a_2 _3809_ (.A1(net84),
    .A2(_0793_),
    .B1(_0888_),
    .B2(_0889_),
    .C1(_0857_),
    .X(net173));
 sky130_fd_sc_hd__a21oi_1 _3810_ (.A1(\core_0.fetch.prev_request_pc[4] ),
    .A2(_0847_),
    .B1(\core_0.fetch.prev_request_pc[5] ),
    .Y(_0890_));
 sky130_fd_sc_hd__nor3_1 _3811_ (.A(_0845_),
    .B(_0848_),
    .C(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__a21o_1 _3812_ (.A1(_0772_),
    .A2(_0861_),
    .B1(_0843_),
    .X(_0892_));
 sky130_fd_sc_hd__o221a_2 _3813_ (.A1(net83),
    .A2(_0793_),
    .B1(_0891_),
    .B2(_0892_),
    .C1(_0857_),
    .X(net172));
 sky130_fd_sc_hd__xnor2_1 _3814_ (.A(\core_0.fetch.prev_request_pc[4] ),
    .B(_0847_),
    .Y(_0893_));
 sky130_fd_sc_hd__nor2_1 _3815_ (.A(_0845_),
    .B(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__a21o_1 _3816_ (.A1(_0763_),
    .A2(_0861_),
    .B1(_0843_),
    .X(_0895_));
 sky130_fd_sc_hd__o221a_2 _3817_ (.A1(net82),
    .A2(_0793_),
    .B1(_0894_),
    .B2(_0895_),
    .C1(_0857_),
    .X(net171));
 sky130_fd_sc_hd__or2_1 _3818_ (.A(\core_0.fetch.prev_request_pc[3] ),
    .B(_0846_),
    .X(_0896_));
 sky130_fd_sc_hd__nor3b_1 _3819_ (.A(_0861_),
    .B(_0847_),
    .C_N(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__a21o_1 _3820_ (.A1(_0761_),
    .A2(_0842_),
    .B1(_0843_),
    .X(_0898_));
 sky130_fd_sc_hd__o221a_2 _3821_ (.A1(net81),
    .A2(_0792_),
    .B1(_0897_),
    .B2(_0898_),
    .C1(_0857_),
    .X(net170));
 sky130_fd_sc_hd__a21oi_1 _3822_ (.A1(\core_0.fetch.prev_request_pc[1] ),
    .A2(\core_0.fetch.prev_request_pc[0] ),
    .B1(\core_0.fetch.prev_request_pc[2] ),
    .Y(_0899_));
 sky130_fd_sc_hd__nor3_1 _3823_ (.A(_0861_),
    .B(_0846_),
    .C(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__a21o_1 _3824_ (.A1(_0766_),
    .A2(_0842_),
    .B1(_0843_),
    .X(_0901_));
 sky130_fd_sc_hd__o221a_4 _3825_ (.A1(net80),
    .A2(_0792_),
    .B1(_0900_),
    .B2(_0901_),
    .C1(_0857_),
    .X(net169));
 sky130_fd_sc_hd__xor2_1 _3826_ (.A(\core_0.fetch.prev_request_pc[1] ),
    .B(\core_0.fetch.prev_request_pc[0] ),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_1 _3827_ (.A0(_0902_),
    .A1(_0759_),
    .S(_0842_),
    .X(_0903_));
 sky130_fd_sc_hd__or2_1 _3828_ (.A(net79),
    .B(_0792_),
    .X(_0904_));
 sky130_fd_sc_hd__o211a_4 _3829_ (.A1(_0862_),
    .A2(_0903_),
    .B1(_0904_),
    .C1(_0858_),
    .X(net168));
 sky130_fd_sc_hd__nor2_1 _3830_ (.A(\core_0.fetch.prev_request_pc[0] ),
    .B(_0845_),
    .Y(_0905_));
 sky130_fd_sc_hd__a21o_1 _3831_ (.A1(_0771_),
    .A2(_0842_),
    .B1(_0843_),
    .X(_0906_));
 sky130_fd_sc_hd__o221a_4 _3832_ (.A1(net72),
    .A2(_0792_),
    .B1(_0905_),
    .B2(_0906_),
    .C1(_0857_),
    .X(net161));
 sky130_fd_sc_hd__inv_2 _3833_ (.A(_0689_),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _3834_ (.A(_0687_),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _3835_ (.A(_0676_),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _3836_ (.A(_0678_),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _3837_ (.A(_0682_),
    .Y(net112));
 sky130_fd_sc_hd__inv_2 _3838_ (.A(_0685_),
    .Y(net113));
 sky130_fd_sc_hd__inv_2 _3839_ (.A(_0681_),
    .Y(net114));
 sky130_fd_sc_hd__inv_2 _3840_ (.A(_0677_),
    .Y(net115));
 sky130_fd_sc_hd__buf_8 _3841_ (.A(net71),
    .X(_0907_));
 sky130_fd_sc_hd__nor2_1 _3842_ (.A(\core_0.decode.input_valid ),
    .B(\core_0.decode.i_submit ),
    .Y(_0908_));
 sky130_fd_sc_hd__nor3_4 _3843_ (.A(_0791_),
    .B(_0747_),
    .C(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__nor2_4 _3844_ (.A(_0907_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__buf_4 _3845_ (.A(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__or3_2 _3846_ (.A(_0791_),
    .B(_0747_),
    .C(_0908_),
    .X(_0912_));
 sky130_fd_sc_hd__nor2_4 _3847_ (.A(net71),
    .B(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__buf_4 _3848_ (.A(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__buf_4 _3849_ (.A(_0914_),
    .X(_0015_));
 sky130_fd_sc_hd__clkinv_2 _3850_ (.A(\core_0.decode.i_instr_l[1] ),
    .Y(_0915_));
 sky130_fd_sc_hd__nor2_1 _3851_ (.A(_0915_),
    .B(\core_0.decode.i_instr_l[0] ),
    .Y(_0916_));
 sky130_fd_sc_hd__or3b_4 _3852_ (.A(\core_0.decode.i_instr_l[6] ),
    .B(\core_0.decode.i_instr_l[5] ),
    .C_N(\core_0.decode.i_instr_l[4] ),
    .X(_0917_));
 sky130_fd_sc_hd__clkbuf_4 _3853_ (.A(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__nand2b_2 _3854_ (.A_N(\core_0.decode.i_instr_l[2] ),
    .B(\core_0.decode.i_instr_l[3] ),
    .Y(_0919_));
 sky130_fd_sc_hd__nor2_1 _3855_ (.A(_0918_),
    .B(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__or3b_1 _3856_ (.A(\core_0.decode.i_instr_l[6] ),
    .B(\core_0.decode.i_instr_l[4] ),
    .C_N(\core_0.decode.i_instr_l[5] ),
    .X(_0921_));
 sky130_fd_sc_hd__clkbuf_4 _3857_ (.A(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__nor2_1 _3858_ (.A(\core_0.decode.i_instr_l[1] ),
    .B(\core_0.decode.i_instr_l[0] ),
    .Y(_0923_));
 sky130_fd_sc_hd__nor2b_2 _3859_ (.A(\core_0.decode.i_instr_l[3] ),
    .B_N(\core_0.decode.i_instr_l[2] ),
    .Y(_0924_));
 sky130_fd_sc_hd__nand2_1 _3860_ (.A(_0923_),
    .B(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__nor2_1 _3861_ (.A(_0922_),
    .B(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__a21o_1 _3862_ (.A1(_0916_),
    .A2(_0920_),
    .B1(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__a22o_1 _3863_ (.A1(\core_0.decode.oc_alu_mode[1] ),
    .A2(_0911_),
    .B1(_0015_),
    .B2(_0927_),
    .X(_0004_));
 sky130_fd_sc_hd__clkbuf_4 _3864_ (.A(\core_0.decode.oc_alu_mode[6] ),
    .X(_0928_));
 sky130_fd_sc_hd__inv_2 _3865_ (.A(\core_0.decode.i_instr_l[0] ),
    .Y(_0929_));
 sky130_fd_sc_hd__nor2_2 _3866_ (.A(\core_0.decode.i_instr_l[1] ),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand2_1 _3867_ (.A(_0924_),
    .B(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__or3_2 _3868_ (.A(\core_0.decode.i_instr_l[1] ),
    .B(\core_0.decode.i_instr_l[0] ),
    .C(_0919_),
    .X(_0932_));
 sky130_fd_sc_hd__a21oi_1 _3869_ (.A1(_0931_),
    .A2(_0932_),
    .B1(_0918_),
    .Y(_0933_));
 sky130_fd_sc_hd__a22o_1 _3870_ (.A1(_0928_),
    .A2(_0911_),
    .B1(_0015_),
    .B2(_0933_),
    .X(_0009_));
 sky130_fd_sc_hd__clkbuf_4 _3871_ (.A(\core_0.decode.oc_alu_mode[7] ),
    .X(_0934_));
 sky130_fd_sc_hd__nor3_4 _3872_ (.A(\core_0.decode.i_instr_l[6] ),
    .B(\core_0.decode.i_instr_l[4] ),
    .C(\core_0.decode.i_instr_l[5] ),
    .Y(_0935_));
 sky130_fd_sc_hd__and2_1 _3873_ (.A(\core_0.decode.i_instr_l[3] ),
    .B(\core_0.decode.i_instr_l[2] ),
    .X(_0936_));
 sky130_fd_sc_hd__and3_1 _3874_ (.A(_0916_),
    .B(_0935_),
    .C(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__nand2_1 _3875_ (.A(\core_0.decode.i_instr_l[1] ),
    .B(_0929_),
    .Y(_0938_));
 sky130_fd_sc_hd__or3_2 _3876_ (.A(\core_0.decode.i_instr_l[3] ),
    .B(\core_0.decode.i_instr_l[2] ),
    .C(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__nand2_1 _3877_ (.A(\core_0.decode.i_instr_l[3] ),
    .B(\core_0.decode.i_instr_l[2] ),
    .Y(_0940_));
 sky130_fd_sc_hd__or3_1 _3878_ (.A(_0915_),
    .B(_0929_),
    .C(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__or3_1 _3879_ (.A(\core_0.decode.i_instr_l[6] ),
    .B(\core_0.decode.i_instr_l[4] ),
    .C(\core_0.decode.i_instr_l[5] ),
    .X(_0942_));
 sky130_fd_sc_hd__buf_2 _3880_ (.A(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__a31o_1 _3881_ (.A1(_0925_),
    .A2(_0939_),
    .A3(_0941_),
    .B1(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__or2b_1 _3882_ (.A(_0937_),
    .B_N(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__nor2_1 _3883_ (.A(\core_0.decode.i_instr_l[3] ),
    .B(\core_0.decode.i_instr_l[2] ),
    .Y(_0946_));
 sky130_fd_sc_hd__nand2_1 _3884_ (.A(_0930_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__nor2_1 _3885_ (.A(_0922_),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__a31o_1 _3886_ (.A1(_0924_),
    .A2(_0930_),
    .A3(_0935_),
    .B1(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__nor2_1 _3887_ (.A(_0917_),
    .B(_0941_),
    .Y(_0950_));
 sky130_fd_sc_hd__or3_1 _3888_ (.A(_0945_),
    .B(_0949_),
    .C(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__a22o_1 _3889_ (.A1(_0934_),
    .A2(_0911_),
    .B1(_0015_),
    .B2(_0951_),
    .X(_0010_));
 sky130_fd_sc_hd__clkbuf_4 _3890_ (.A(_0913_),
    .X(_0952_));
 sky130_fd_sc_hd__and3b_1 _3891_ (.A_N(_0917_),
    .B(_0936_),
    .C(_0915_),
    .X(_0953_));
 sky130_fd_sc_hd__clkbuf_4 _3892_ (.A(_0910_),
    .X(_0954_));
 sky130_fd_sc_hd__buf_4 _3893_ (.A(\core_0.execute.alu_mul_div.i_mul ),
    .X(_0955_));
 sky130_fd_sc_hd__a32o_1 _3894_ (.A1(_0929_),
    .A2(_0952_),
    .A3(_0953_),
    .B1(_0954_),
    .B2(_0955_),
    .X(_0011_));
 sky130_fd_sc_hd__clkbuf_4 _3895_ (.A(\core_0.decode.oc_alu_mode[9] ),
    .X(_0956_));
 sky130_fd_sc_hd__and3_1 _3896_ (.A(\core_0.decode.i_instr_l[1] ),
    .B(\core_0.decode.i_instr_l[0] ),
    .C(_0924_),
    .X(_0957_));
 sky130_fd_sc_hd__or2b_1 _3897_ (.A(_0917_),
    .B_N(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__o21ai_1 _3898_ (.A1(_0925_),
    .A2(_0918_),
    .B1(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__a22o_1 _3899_ (.A1(_0956_),
    .A2(_0911_),
    .B1(_0015_),
    .B2(_0959_),
    .X(_0012_));
 sky130_fd_sc_hd__buf_4 _3900_ (.A(\core_0.execute.alu_mul_div.i_mod ),
    .X(_0960_));
 sky130_fd_sc_hd__and3b_1 _3901_ (.A_N(_0922_),
    .B(_0923_),
    .C(_0936_),
    .X(_0961_));
 sky130_fd_sc_hd__a22o_1 _3902_ (.A1(_0960_),
    .A2(_0911_),
    .B1(_0015_),
    .B2(_0961_),
    .X(_0000_));
 sky130_fd_sc_hd__clkbuf_4 _3903_ (.A(\core_0.decode.oc_alu_mode[4] ),
    .X(_0962_));
 sky130_fd_sc_hd__or3b_1 _3904_ (.A(_0915_),
    .B(_0929_),
    .C_N(_0946_),
    .X(_0963_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3905_ (.A(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__a21oi_1 _3906_ (.A1(_0932_),
    .A2(_0964_),
    .B1(_0943_),
    .Y(_0965_));
 sky130_fd_sc_hd__nor3_1 _3907_ (.A(_0929_),
    .B(_0919_),
    .C(_0943_),
    .Y(_0966_));
 sky130_fd_sc_hd__and2_1 _3908_ (.A(_0915_),
    .B(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__and2_1 _3909_ (.A(_0935_),
    .B(_0957_),
    .X(_0968_));
 sky130_fd_sc_hd__or2_1 _3910_ (.A(_0967_),
    .B(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__or2_1 _3911_ (.A(_0965_),
    .B(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__nor2_1 _3912_ (.A(_0922_),
    .B(_0939_),
    .Y(_0971_));
 sky130_fd_sc_hd__nand2_1 _3913_ (.A(_0924_),
    .B(_0916_),
    .Y(_0972_));
 sky130_fd_sc_hd__nor2_1 _3914_ (.A(_0943_),
    .B(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__or2_1 _3915_ (.A(_0971_),
    .B(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__and3b_1 _3916_ (.A_N(_0922_),
    .B(_0923_),
    .C(_0946_),
    .X(_0975_));
 sky130_fd_sc_hd__nor2_2 _3917_ (.A(_0922_),
    .B(_0919_),
    .Y(_0976_));
 sky130_fd_sc_hd__or4_1 _3918_ (.A(_0970_),
    .B(_0974_),
    .C(_0975_),
    .D(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__a22o_1 _3919_ (.A1(_0962_),
    .A2(_0911_),
    .B1(_0015_),
    .B2(_0977_),
    .X(_0007_));
 sky130_fd_sc_hd__buf_4 _3920_ (.A(\core_0.decode.oc_alu_mode[11] ),
    .X(_0978_));
 sky130_fd_sc_hd__and3_1 _3921_ (.A(_0930_),
    .B(_0935_),
    .C(_0936_),
    .X(_0979_));
 sky130_fd_sc_hd__a21o_1 _3922_ (.A1(\core_0.decode.i_instr_l[1] ),
    .A2(_0966_),
    .B1(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__nor3_1 _3923_ (.A(_0938_),
    .B(_0919_),
    .C(_0943_),
    .Y(_0981_));
 sky130_fd_sc_hd__a31o_1 _3924_ (.A1(_0923_),
    .A2(_0935_),
    .A3(_0936_),
    .B1(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__or2_1 _3925_ (.A(_0980_),
    .B(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__a22o_1 _3926_ (.A1(_0978_),
    .A2(_0911_),
    .B1(_0015_),
    .B2(_0983_),
    .X(_0001_));
 sky130_fd_sc_hd__buf_4 _3927_ (.A(\core_0.decode.oc_alu_mode[12] ),
    .X(_0984_));
 sky130_fd_sc_hd__nor2_1 _3928_ (.A(_0922_),
    .B(_0931_),
    .Y(_0985_));
 sky130_fd_sc_hd__nor2_1 _3929_ (.A(_0922_),
    .B(_0972_),
    .Y(_0986_));
 sky130_fd_sc_hd__or2_1 _3930_ (.A(_0985_),
    .B(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__a22o_1 _3931_ (.A1(_0984_),
    .A2(_0911_),
    .B1(_0015_),
    .B2(_0987_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_4 _3932_ (.A(\core_0.execute.alu_mul_div.i_div ),
    .X(_0988_));
 sky130_fd_sc_hd__buf_4 _3933_ (.A(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__a32o_1 _3934_ (.A1(\core_0.decode.i_instr_l[0] ),
    .A2(_0952_),
    .A3(_0953_),
    .B1(_0954_),
    .B2(_0989_),
    .X(_0008_));
 sky130_fd_sc_hd__buf_4 _3935_ (.A(_0910_),
    .X(_0990_));
 sky130_fd_sc_hd__nor2_1 _3936_ (.A(_0922_),
    .B(_0964_),
    .Y(_0991_));
 sky130_fd_sc_hd__a21o_1 _3937_ (.A1(_0920_),
    .A2(_0930_),
    .B1(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__a22o_1 _3938_ (.A1(\core_0.decode.oc_alu_mode[13] ),
    .A2(_0990_),
    .B1(_0015_),
    .B2(_0992_),
    .X(_0003_));
 sky130_fd_sc_hd__or2b_1 _3939_ (.A(_0922_),
    .B_N(_0957_),
    .X(_0993_));
 sky130_fd_sc_hd__nand2_1 _3940_ (.A(_0909_),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__buf_4 _3941_ (.A(_0665_),
    .X(_0995_));
 sky130_fd_sc_hd__buf_6 _3942_ (.A(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__buf_6 _3943_ (.A(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__o211a_1 _3944_ (.A1(\core_0.decode.oc_alu_mode[3] ),
    .A2(_0909_),
    .B1(_0994_),
    .C1(_0997_),
    .X(_0006_));
 sky130_fd_sc_hd__clkbuf_4 _3945_ (.A(\core_0.decode.oc_alu_mode[2] ),
    .X(_0998_));
 sky130_fd_sc_hd__buf_4 _3946_ (.A(_0914_),
    .X(_0999_));
 sky130_fd_sc_hd__nor2_1 _3947_ (.A(_0918_),
    .B(_0972_),
    .Y(_1000_));
 sky130_fd_sc_hd__and3_1 _3948_ (.A(\core_0.decode.i_instr_l[1] ),
    .B(\core_0.decode.i_instr_l[0] ),
    .C(_0920_),
    .X(_1001_));
 sky130_fd_sc_hd__nor2_1 _3949_ (.A(_0918_),
    .B(_0964_),
    .Y(_1002_));
 sky130_fd_sc_hd__or3_1 _3950_ (.A(_1000_),
    .B(_1001_),
    .C(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__a22o_1 _3951_ (.A1(_0998_),
    .A2(_0990_),
    .B1(_0999_),
    .B2(_1003_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _3952_ (.A0(\core_0.fetch.prev_req_branch_pred ),
    .A1(_0841_),
    .S(net70),
    .X(_1004_));
 sky130_fd_sc_hd__clkbuf_1 _3953_ (.A(_1004_),
    .X(\core_0.fetch.current_req_branch_pred ));
 sky130_fd_sc_hd__nand2_4 _3954_ (.A(\core_0.ew_addr[0] ),
    .B(\core_0.ew_mem_width ),
    .Y(_1005_));
 sky130_fd_sc_hd__clkbuf_4 _3955_ (.A(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__clkbuf_4 _3956_ (.A(_1006_),
    .X(net157));
 sky130_fd_sc_hd__and2_1 _3957_ (.A(\core_0.ew_data[0] ),
    .B(net157),
    .X(_1007_));
 sky130_fd_sc_hd__clkbuf_1 _3958_ (.A(_1007_),
    .X(net139));
 sky130_fd_sc_hd__and2_1 _3959_ (.A(\core_0.ew_data[1] ),
    .B(net157),
    .X(_1008_));
 sky130_fd_sc_hd__clkbuf_1 _3960_ (.A(_1008_),
    .X(net146));
 sky130_fd_sc_hd__and2_1 _3961_ (.A(\core_0.ew_data[2] ),
    .B(net157),
    .X(_1009_));
 sky130_fd_sc_hd__clkbuf_1 _3962_ (.A(_1009_),
    .X(net147));
 sky130_fd_sc_hd__and2_1 _3963_ (.A(\core_0.ew_data[3] ),
    .B(net157),
    .X(_1010_));
 sky130_fd_sc_hd__clkbuf_1 _3964_ (.A(_1010_),
    .X(net148));
 sky130_fd_sc_hd__and2_1 _3965_ (.A(\core_0.ew_data[4] ),
    .B(net157),
    .X(_1011_));
 sky130_fd_sc_hd__clkbuf_1 _3966_ (.A(_1011_),
    .X(net149));
 sky130_fd_sc_hd__and2_1 _3967_ (.A(\core_0.ew_data[5] ),
    .B(net157),
    .X(_1012_));
 sky130_fd_sc_hd__clkbuf_1 _3968_ (.A(_1012_),
    .X(net150));
 sky130_fd_sc_hd__and2_1 _3969_ (.A(\core_0.ew_data[6] ),
    .B(net157),
    .X(_1013_));
 sky130_fd_sc_hd__clkbuf_1 _3970_ (.A(_1013_),
    .X(net151));
 sky130_fd_sc_hd__and2_1 _3971_ (.A(\core_0.ew_data[7] ),
    .B(net157),
    .X(_1014_));
 sky130_fd_sc_hd__clkbuf_1 _3972_ (.A(_1014_),
    .X(net152));
 sky130_fd_sc_hd__mux2_1 _3973_ (.A0(\core_0.ew_data[0] ),
    .A1(\core_0.ew_data[8] ),
    .S(net157),
    .X(_1015_));
 sky130_fd_sc_hd__clkbuf_1 _3974_ (.A(_1015_),
    .X(net153));
 sky130_fd_sc_hd__mux2_1 _3975_ (.A0(\core_0.ew_data[1] ),
    .A1(\core_0.ew_data[9] ),
    .S(_1006_),
    .X(_1016_));
 sky130_fd_sc_hd__clkbuf_1 _3976_ (.A(_1016_),
    .X(net154));
 sky130_fd_sc_hd__mux2_1 _3977_ (.A0(\core_0.ew_data[2] ),
    .A1(\core_0.ew_data[10] ),
    .S(_1006_),
    .X(_1017_));
 sky130_fd_sc_hd__clkbuf_1 _3978_ (.A(_1017_),
    .X(net140));
 sky130_fd_sc_hd__mux2_1 _3979_ (.A0(\core_0.ew_data[3] ),
    .A1(\core_0.ew_data[11] ),
    .S(_1006_),
    .X(_1018_));
 sky130_fd_sc_hd__clkbuf_1 _3980_ (.A(_1018_),
    .X(net141));
 sky130_fd_sc_hd__mux2_1 _3981_ (.A0(\core_0.ew_data[4] ),
    .A1(\core_0.ew_data[12] ),
    .S(_1006_),
    .X(_1019_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3982_ (.A(_1019_),
    .X(net142));
 sky130_fd_sc_hd__mux2_1 _3983_ (.A0(\core_0.ew_data[5] ),
    .A1(\core_0.ew_data[13] ),
    .S(_1006_),
    .X(_1020_));
 sky130_fd_sc_hd__clkbuf_1 _3984_ (.A(_1020_),
    .X(net143));
 sky130_fd_sc_hd__mux2_2 _3985_ (.A0(\core_0.ew_data[6] ),
    .A1(\core_0.ew_data[14] ),
    .S(_1006_),
    .X(_1021_));
 sky130_fd_sc_hd__clkbuf_1 _3986_ (.A(_1021_),
    .X(net144));
 sky130_fd_sc_hd__mux2_2 _3987_ (.A0(\core_0.ew_data[7] ),
    .A1(\core_0.ew_data[15] ),
    .S(_1006_),
    .X(_1022_));
 sky130_fd_sc_hd__clkbuf_1 _3988_ (.A(_1022_),
    .X(net145));
 sky130_fd_sc_hd__or2b_2 _3989_ (.A(\core_0.ew_addr[0] ),
    .B_N(\core_0.ew_mem_width ),
    .X(_1023_));
 sky130_fd_sc_hd__clkbuf_1 _3990_ (.A(_1023_),
    .X(net158));
 sky130_fd_sc_hd__inv_2 _3991_ (.A(net17),
    .Y(net160));
 sky130_fd_sc_hd__nor2_2 _3992_ (.A(_0791_),
    .B(\core_0.fetch.flush_event_invalidate ),
    .Y(_1024_));
 sky130_fd_sc_hd__o211ai_4 _3993_ (.A1(_0670_),
    .A2(net70),
    .B1(_0748_),
    .C1(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__inv_2 _3994_ (.A(_1025_),
    .Y(\core_0.fetch.submitable ));
 sky130_fd_sc_hd__and2_2 _3995_ (.A(net155),
    .B(\core_0.ew_addr_high[0] ),
    .X(_1026_));
 sky130_fd_sc_hd__clkbuf_1 _3996_ (.A(_1026_),
    .X(net122));
 sky130_fd_sc_hd__buf_6 _3997_ (.A(_0746_),
    .X(_1027_));
 sky130_fd_sc_hd__buf_4 _3998_ (.A(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__inv_2 _3999_ (.A(\core_0.execute.sreg_jtr_buff.o_d[0] ),
    .Y(_1029_));
 sky130_fd_sc_hd__nor3_4 _4000_ (.A(net181),
    .B(net184),
    .C(net183),
    .Y(_1030_));
 sky130_fd_sc_hd__nor4_4 _4001_ (.A(net193),
    .B(net180),
    .C(net179),
    .D(net182),
    .Y(_1031_));
 sky130_fd_sc_hd__and4bb_1 _4002_ (.A_N(net185),
    .B_N(net192),
    .C(_1030_),
    .D(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__clkbuf_2 _4003_ (.A(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__nor4_4 _4004_ (.A(net189),
    .B(net188),
    .C(net191),
    .D(net190),
    .Y(_1034_));
 sky130_fd_sc_hd__and2b_1 _4005_ (.A_N(net178),
    .B(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__nor2_1 _4006_ (.A(net187),
    .B(net186),
    .Y(_1036_));
 sky130_fd_sc_hd__and3_2 _4007_ (.A(_1033_),
    .B(_1035_),
    .C(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__buf_4 _4008_ (.A(\core_0.dec_sreg_irt ),
    .X(_1038_));
 sky130_fd_sc_hd__a21o_2 _4009_ (.A1(\core_0.dec_sreg_store ),
    .A2(_1037_),
    .B1(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__o21a_4 _4010_ (.A1(\core_0.dec_jump_cond_code[4] ),
    .A2(_1039_),
    .B1(_0746_),
    .X(_1040_));
 sky130_fd_sc_hd__and4_1 _4011_ (.A(\core_0.dec_sreg_store ),
    .B(_1030_),
    .C(_1031_),
    .D(_1034_),
    .X(_1041_));
 sky130_fd_sc_hd__and3_1 _4012_ (.A(net192),
    .B(_0746_),
    .C(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__a211o_1 _4013_ (.A1(_1029_),
    .A2(_1040_),
    .B1(_1042_),
    .C1(_0674_),
    .X(_1043_));
 sky130_fd_sc_hd__and3b_1 _4014_ (.A_N(net106),
    .B(\core_0.execute.sreg_jtr_buff.o_d[0] ),
    .C(_1040_),
    .X(_1044_));
 sky130_fd_sc_hd__a211o_1 _4015_ (.A1(net106),
    .A2(_1043_),
    .B1(_1044_),
    .C1(_0693_),
    .X(_1045_));
 sky130_fd_sc_hd__inv_2 _4016_ (.A(\core_0.execute.alu_flag_reg.o_d[2] ),
    .Y(_1046_));
 sky130_fd_sc_hd__xor2_1 _4017_ (.A(\core_0.dec_jump_cond_code[1] ),
    .B(\core_0.dec_jump_cond_code[0] ),
    .X(_1047_));
 sky130_fd_sc_hd__inv_2 _4018_ (.A(\core_0.execute.alu_flag_reg.o_d[0] ),
    .Y(_1048_));
 sky130_fd_sc_hd__o221a_1 _4019_ (.A1(_1046_),
    .A2(\core_0.dec_jump_cond_code[0] ),
    .B1(_1047_),
    .B2(_1048_),
    .C1(\core_0.dec_jump_cond_code[2] ),
    .X(_1049_));
 sky130_fd_sc_hd__inv_2 _4020_ (.A(\core_0.dec_jump_cond_code[0] ),
    .Y(_1050_));
 sky130_fd_sc_hd__or4_1 _4021_ (.A(\core_0.execute.alu_flag_reg.o_d[2] ),
    .B(\core_0.execute.alu_flag_reg.o_d[0] ),
    .C(\core_0.dec_jump_cond_code[1] ),
    .D(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__a31o_1 _4022_ (.A1(_1048_),
    .A2(\core_0.dec_jump_cond_code[1] ),
    .A3(_1050_),
    .B1(\core_0.dec_jump_cond_code[2] ),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_1 _4023_ (.A0(\core_0.execute.alu_flag_reg.o_d[1] ),
    .A1(\core_0.execute.alu_flag_reg.o_d[2] ),
    .S(\core_0.dec_jump_cond_code[1] ),
    .X(_1053_));
 sky130_fd_sc_hd__nor2_1 _4024_ (.A(_1050_),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__o2bb2a_1 _4025_ (.A1_N(_1049_),
    .A2_N(_1051_),
    .B1(_1052_),
    .B2(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__a21o_1 _4026_ (.A1(\core_0.execute.alu_flag_reg.o_d[0] ),
    .A2(_1050_),
    .B1(\core_0.execute.alu_flag_reg.o_d[1] ),
    .X(_1056_));
 sky130_fd_sc_hd__or4_1 _4027_ (.A(\core_0.execute.alu_flag_reg.o_d[3] ),
    .B(\core_0.dec_jump_cond_code[2] ),
    .C(\core_0.dec_jump_cond_code[1] ),
    .D(\core_0.dec_jump_cond_code[0] ),
    .X(_1057_));
 sky130_fd_sc_hd__o31ai_1 _4028_ (.A1(\core_0.execute.alu_flag_reg.o_d[4] ),
    .A2(\core_0.dec_jump_cond_code[1] ),
    .A3(_1050_),
    .B1(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__nor2_1 _4029_ (.A(\core_0.execute.alu_flag_reg.o_d[1] ),
    .B(\core_0.execute.alu_flag_reg.o_d[0] ),
    .Y(_1059_));
 sky130_fd_sc_hd__o21a_1 _4030_ (.A1(\core_0.dec_jump_cond_code[0] ),
    .A2(_1059_),
    .B1(\core_0.dec_jump_cond_code[2] ),
    .X(_1060_));
 sky130_fd_sc_hd__a211o_1 _4031_ (.A1(\core_0.dec_jump_cond_code[1] ),
    .A2(_1056_),
    .B1(_1058_),
    .C1(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__mux2_2 _4032_ (.A0(_1055_),
    .A1(_1061_),
    .S(\core_0.dec_jump_cond_code[3] ),
    .X(_1062_));
 sky130_fd_sc_hd__a31o_1 _4033_ (.A1(\core_0.dec_jump_cond_code[4] ),
    .A2(\core_0.de_jmp_pred ),
    .A3(_1062_),
    .B1(_1039_),
    .X(_1063_));
 sky130_fd_sc_hd__or3b_1 _4034_ (.A(\core_0.de_jmp_pred ),
    .B(_1062_),
    .C_N(\core_0.dec_jump_cond_code[4] ),
    .X(_1064_));
 sky130_fd_sc_hd__or3b_1 _4035_ (.A(_1045_),
    .B(_1063_),
    .C_N(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__a21o_1 _4036_ (.A1(_1028_),
    .A2(_1065_),
    .B1(_0694_),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_4 _4037_ (.A(_0995_),
    .X(_1066_));
 sky130_fd_sc_hd__and2_1 _4038_ (.A(_1066_),
    .B(_1045_),
    .X(_1067_));
 sky130_fd_sc_hd__clkbuf_1 _4039_ (.A(_1067_),
    .X(_0014_));
 sky130_fd_sc_hd__or3_1 _4040_ (.A(_0791_),
    .B(_0694_),
    .C(_0695_),
    .X(_1068_));
 sky130_fd_sc_hd__buf_4 _4041_ (.A(_0738_),
    .X(_1069_));
 sky130_fd_sc_hd__buf_4 _4042_ (.A(_0745_),
    .X(_1070_));
 sky130_fd_sc_hd__nor3_4 _4043_ (.A(_1068_),
    .B(_1069_),
    .C(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__and3_1 _4044_ (.A(\core_0.execute.sreg_priv_control.o_d[0] ),
    .B(\core_0.dec_sreg_store ),
    .C(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__clkbuf_1 _4045_ (.A(_1072_),
    .X(net210));
 sky130_fd_sc_hd__or4_2 _4046_ (.A(_0912_),
    .B(_0938_),
    .C(_0918_),
    .D(_0940_),
    .X(_1073_));
 sky130_fd_sc_hd__or4_1 _4047_ (.A(_0915_),
    .B(_0912_),
    .C(_0943_),
    .D(_0940_),
    .X(_1074_));
 sky130_fd_sc_hd__buf_6 _4048_ (.A(_0995_),
    .X(_1075_));
 sky130_fd_sc_hd__o2111a_1 _4049_ (.A1(\core_0.dec_pc_inc ),
    .A2(_0909_),
    .B1(_1073_),
    .C1(_1074_),
    .D1(_1075_),
    .X(_0016_));
 sky130_fd_sc_hd__buf_4 _4050_ (.A(\core_0.dec_r_bus_imm ),
    .X(_1076_));
 sky130_fd_sc_hd__buf_6 _4051_ (.A(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__nor2_1 _4052_ (.A(_0932_),
    .B(_0943_),
    .Y(_1078_));
 sky130_fd_sc_hd__o21ai_1 _4053_ (.A1(_0917_),
    .A2(_0932_),
    .B1(_0958_),
    .Y(_1079_));
 sky130_fd_sc_hd__or4_1 _4054_ (.A(_1078_),
    .B(_0973_),
    .C(_0976_),
    .D(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__or4_1 _4055_ (.A(_0980_),
    .B(_1000_),
    .C(_1001_),
    .D(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__or2_1 _4056_ (.A(_0926_),
    .B(_0991_),
    .X(_1082_));
 sky130_fd_sc_hd__or3_1 _4057_ (.A(_0986_),
    .B(_1001_),
    .C(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__or2_1 _4058_ (.A(_0950_),
    .B(_0975_),
    .X(_1084_));
 sky130_fd_sc_hd__or3_1 _4059_ (.A(_0948_),
    .B(_0971_),
    .C(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__a41o_1 _4060_ (.A1(_0931_),
    .A2(_0939_),
    .A3(_0964_),
    .A4(_0972_),
    .B1(_0943_),
    .X(_1086_));
 sky130_fd_sc_hd__or2b_1 _4061_ (.A(_1085_),
    .B_N(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__or4_1 _4062_ (.A(_0945_),
    .B(_1081_),
    .C(_1083_),
    .D(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__a22o_1 _4063_ (.A1(_1077_),
    .A2(_0990_),
    .B1(_0999_),
    .B2(_1088_),
    .X(_0017_));
 sky130_fd_sc_hd__o21a_1 _4064_ (.A1(_0916_),
    .A2(_0930_),
    .B1(_0920_),
    .X(_1089_));
 sky130_fd_sc_hd__or3_1 _4065_ (.A(_0991_),
    .B(_1001_),
    .C(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__or3b_1 _4066_ (.A(_0987_),
    .B(_1082_),
    .C_N(_0993_),
    .X(_1091_));
 sky130_fd_sc_hd__nor2_1 _4067_ (.A(_0918_),
    .B(_0931_),
    .Y(_1092_));
 sky130_fd_sc_hd__or3_1 _4068_ (.A(_1092_),
    .B(_1000_),
    .C(_1079_),
    .X(_1093_));
 sky130_fd_sc_hd__a21oi_1 _4069_ (.A1(_0925_),
    .A2(_0964_),
    .B1(_0918_),
    .Y(_1094_));
 sky130_fd_sc_hd__or4_1 _4070_ (.A(_1078_),
    .B(_0969_),
    .C(_1093_),
    .D(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__or4_1 _4071_ (.A(_0983_),
    .B(_1090_),
    .C(_1091_),
    .D(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__a22o_1 _4072_ (.A1(\core_0.dec_alu_flags_ie ),
    .A2(_0990_),
    .B1(_0999_),
    .B2(_1096_),
    .X(_0018_));
 sky130_fd_sc_hd__a22o_1 _4073_ (.A1(\core_0.dec_alu_carry_en ),
    .A2(_0990_),
    .B1(_0999_),
    .B2(_0966_),
    .X(_0019_));
 sky130_fd_sc_hd__a21o_2 _4074_ (.A1(\core_0.decode.i_instr_l[0] ),
    .A2(_0976_),
    .B1(_0974_),
    .X(_1097_));
 sky130_fd_sc_hd__or3_1 _4075_ (.A(_0953_),
    .B(_1079_),
    .C(_1090_),
    .X(_1098_));
 sky130_fd_sc_hd__inv_2 _4076_ (.A(_0947_),
    .Y(_1099_));
 sky130_fd_sc_hd__a221o_1 _4077_ (.A1(_0935_),
    .A2(_1099_),
    .B1(_0976_),
    .B2(_0929_),
    .C1(_0975_),
    .X(_1100_));
 sky130_fd_sc_hd__or4_1 _4078_ (.A(_0961_),
    .B(_0970_),
    .C(_1091_),
    .D(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__or3_4 _4079_ (.A(_1096_),
    .B(_1098_),
    .C(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__a22o_1 _4080_ (.A1(\core_0.decode.i_instr_l[13] ),
    .A2(_1097_),
    .B1(_1102_),
    .B2(\core_0.decode.i_instr_l[10] ),
    .X(_1103_));
 sky130_fd_sc_hd__a22o_1 _4081_ (.A1(_0715_),
    .A2(_0990_),
    .B1(_0999_),
    .B2(_1103_),
    .X(_0020_));
 sky130_fd_sc_hd__a22o_1 _4082_ (.A1(\core_0.decode.i_instr_l[14] ),
    .A2(_1097_),
    .B1(_1102_),
    .B2(\core_0.decode.i_instr_l[11] ),
    .X(_1104_));
 sky130_fd_sc_hd__a22o_1 _4083_ (.A1(_0704_),
    .A2(_0990_),
    .B1(_0999_),
    .B2(_1104_),
    .X(_0021_));
 sky130_fd_sc_hd__a22o_1 _4084_ (.A1(\core_0.decode.i_instr_l[15] ),
    .A2(_1097_),
    .B1(_1102_),
    .B2(\core_0.decode.i_instr_l[12] ),
    .X(_1105_));
 sky130_fd_sc_hd__a22o_1 _4085_ (.A1(_0706_),
    .A2(_0990_),
    .B1(_0999_),
    .B2(_1105_),
    .X(_0022_));
 sky130_fd_sc_hd__nor2_1 _4086_ (.A(_0918_),
    .B(_0947_),
    .Y(_1106_));
 sky130_fd_sc_hd__or2_1 _4087_ (.A(_0949_),
    .B(_1097_),
    .X(_1107_));
 sky130_fd_sc_hd__or2_2 _4088_ (.A(_1106_),
    .B(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__or4_1 _4089_ (.A(_1092_),
    .B(_0953_),
    .C(_0961_),
    .D(_0985_),
    .X(_1109_));
 sky130_fd_sc_hd__or3_1 _4090_ (.A(_1094_),
    .B(_1089_),
    .C(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__or4_4 _4091_ (.A(_0966_),
    .B(_0968_),
    .C(_0982_),
    .D(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__a22o_1 _4092_ (.A1(\core_0.decode.i_instr_l[10] ),
    .A2(_1108_),
    .B1(_1111_),
    .B2(\core_0.decode.i_instr_l[13] ),
    .X(_1112_));
 sky130_fd_sc_hd__a22o_1 _4093_ (.A1(_0571_),
    .A2(_0990_),
    .B1(_0999_),
    .B2(_1112_),
    .X(_0023_));
 sky130_fd_sc_hd__a22o_1 _4094_ (.A1(\core_0.decode.i_instr_l[11] ),
    .A2(_1108_),
    .B1(_1111_),
    .B2(\core_0.decode.i_instr_l[14] ),
    .X(_1113_));
 sky130_fd_sc_hd__a22o_1 _4095_ (.A1(_0569_),
    .A2(_0990_),
    .B1(_0999_),
    .B2(_1113_),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_4 _4096_ (.A(_0910_),
    .X(_1114_));
 sky130_fd_sc_hd__a22o_1 _4097_ (.A1(\core_0.decode.i_instr_l[12] ),
    .A2(_1108_),
    .B1(_1111_),
    .B2(\core_0.decode.i_instr_l[15] ),
    .X(_1115_));
 sky130_fd_sc_hd__a22o_1 _4098_ (.A1(_0573_),
    .A2(_1114_),
    .B1(_0999_),
    .B2(_1115_),
    .X(_0025_));
 sky130_fd_sc_hd__and4b_1 _4099_ (.A_N(_0917_),
    .B(_0946_),
    .C(_0915_),
    .D(_0929_),
    .X(_1116_));
 sky130_fd_sc_hd__or4_1 _4100_ (.A(_0967_),
    .B(_0981_),
    .C(_1084_),
    .D(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__or4b_1 _4101_ (.A(_1093_),
    .B(_1094_),
    .C(_1117_),
    .D_N(_0944_),
    .X(_1118_));
 sky130_fd_sc_hd__or3_2 _4102_ (.A(_1101_),
    .B(_1110_),
    .C(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__and2b_1 _4103_ (.A_N(\core_0.decode.i_instr_l[8] ),
    .B(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__and3b_1 _4104_ (.A_N(\core_0.decode.i_instr_l[7] ),
    .B(_0909_),
    .C(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__buf_6 _4105_ (.A(_0907_),
    .X(_1122_));
 sky130_fd_sc_hd__nor2_2 _4106_ (.A(_1122_),
    .B(\core_0.decode.i_instr_l[9] ),
    .Y(_1123_));
 sky130_fd_sc_hd__a22o_1 _4107_ (.A1(\core_0.dec_rf_ie[0] ),
    .A2(_1114_),
    .B1(_1121_),
    .B2(_1123_),
    .X(_0026_));
 sky130_fd_sc_hd__and3_1 _4108_ (.A(\core_0.decode.i_instr_l[7] ),
    .B(_0909_),
    .C(_1120_),
    .X(_1124_));
 sky130_fd_sc_hd__a22o_1 _4109_ (.A1(\core_0.dec_rf_ie[1] ),
    .A2(_1114_),
    .B1(_1123_),
    .B2(_1124_),
    .X(_0027_));
 sky130_fd_sc_hd__and4b_1 _4110_ (.A_N(\core_0.decode.i_instr_l[7] ),
    .B(_0909_),
    .C(_1119_),
    .D(\core_0.decode.i_instr_l[8] ),
    .X(_1125_));
 sky130_fd_sc_hd__a22o_1 _4111_ (.A1(\core_0.dec_rf_ie[2] ),
    .A2(_1114_),
    .B1(_1123_),
    .B2(_1125_),
    .X(_0028_));
 sky130_fd_sc_hd__and4_1 _4112_ (.A(\core_0.decode.i_instr_l[8] ),
    .B(\core_0.decode.i_instr_l[7] ),
    .C(_0909_),
    .D(_1119_),
    .X(_1126_));
 sky130_fd_sc_hd__a22o_1 _4113_ (.A1(\core_0.dec_rf_ie[3] ),
    .A2(_1114_),
    .B1(_1123_),
    .B2(_1126_),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _4114_ (.A(_0995_),
    .B(\core_0.decode.i_instr_l[9] ),
    .X(_1127_));
 sky130_fd_sc_hd__a22o_1 _4115_ (.A1(\core_0.dec_rf_ie[4] ),
    .A2(_1114_),
    .B1(_1121_),
    .B2(_1127_),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _4116_ (.A1(\core_0.dec_rf_ie[5] ),
    .A2(_1114_),
    .B1(_1124_),
    .B2(_1127_),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_1 _4117_ (.A1(\core_0.dec_rf_ie[6] ),
    .A2(_1114_),
    .B1(_1125_),
    .B2(_1127_),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_1 _4118_ (.A1(\core_0.dec_rf_ie[7] ),
    .A2(_1114_),
    .B1(_1126_),
    .B2(_1127_),
    .X(_0033_));
 sky130_fd_sc_hd__a32o_1 _4119_ (.A1(\core_0.decode.i_instr_l[7] ),
    .A2(_0914_),
    .A3(_0937_),
    .B1(_0954_),
    .B2(\core_0.dec_jump_cond_code[0] ),
    .X(_0034_));
 sky130_fd_sc_hd__a32o_1 _4120_ (.A1(\core_0.decode.i_instr_l[8] ),
    .A2(_0914_),
    .A3(_0937_),
    .B1(_0910_),
    .B2(\core_0.dec_jump_cond_code[1] ),
    .X(_0035_));
 sky130_fd_sc_hd__a32o_1 _4121_ (.A1(\core_0.decode.i_instr_l[9] ),
    .A2(_0914_),
    .A3(_0937_),
    .B1(_0910_),
    .B2(\core_0.dec_jump_cond_code[2] ),
    .X(_0036_));
 sky130_fd_sc_hd__a32o_1 _4122_ (.A1(\core_0.decode.i_instr_l[10] ),
    .A2(_0914_),
    .A3(_0937_),
    .B1(_0910_),
    .B2(\core_0.dec_jump_cond_code[3] ),
    .X(_0037_));
 sky130_fd_sc_hd__buf_4 _4123_ (.A(_1122_),
    .X(_1128_));
 sky130_fd_sc_hd__a2bb2o_1 _4124_ (.A1_N(_1128_),
    .A2_N(_1074_),
    .B1(_0911_),
    .B2(\core_0.dec_jump_cond_code[4] ),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _4125_ (.A0(net178),
    .A1(\core_0.decode.i_imm_pass[0] ),
    .S(_0914_),
    .X(_1129_));
 sky130_fd_sc_hd__clkbuf_1 _4126_ (.A(_1129_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _4127_ (.A0(net185),
    .A1(\core_0.decode.i_imm_pass[1] ),
    .S(_0914_),
    .X(_1130_));
 sky130_fd_sc_hd__clkbuf_1 _4128_ (.A(_1130_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _4129_ (.A0(net186),
    .A1(\core_0.decode.i_imm_pass[2] ),
    .S(_0914_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_1 _4130_ (.A(_1131_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _4131_ (.A0(net187),
    .A1(\core_0.decode.i_imm_pass[3] ),
    .S(_0914_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _4132_ (.A(_1132_),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_4 _4133_ (.A(_0913_),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _4134_ (.A0(net188),
    .A1(\core_0.decode.i_imm_pass[4] ),
    .S(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _4135_ (.A(_1134_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _4136_ (.A0(net189),
    .A1(\core_0.decode.i_imm_pass[5] ),
    .S(_1133_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_1 _4137_ (.A(_1135_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _4138_ (.A0(net190),
    .A1(\core_0.decode.i_imm_pass[6] ),
    .S(_1133_),
    .X(_1136_));
 sky130_fd_sc_hd__clkbuf_1 _4139_ (.A(_1136_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _4140_ (.A0(net191),
    .A1(\core_0.decode.i_imm_pass[7] ),
    .S(_1133_),
    .X(_1137_));
 sky130_fd_sc_hd__clkbuf_1 _4141_ (.A(_1137_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _4142_ (.A0(net192),
    .A1(\core_0.decode.i_imm_pass[8] ),
    .S(_1133_),
    .X(_1138_));
 sky130_fd_sc_hd__clkbuf_1 _4143_ (.A(_1138_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _4144_ (.A0(net193),
    .A1(\core_0.decode.i_imm_pass[9] ),
    .S(_1133_),
    .X(_1139_));
 sky130_fd_sc_hd__clkbuf_1 _4145_ (.A(_1139_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _4146_ (.A0(net179),
    .A1(\core_0.decode.i_imm_pass[10] ),
    .S(_1133_),
    .X(_1140_));
 sky130_fd_sc_hd__clkbuf_1 _4147_ (.A(_1140_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _4148_ (.A0(net180),
    .A1(\core_0.decode.i_imm_pass[11] ),
    .S(_1133_),
    .X(_1141_));
 sky130_fd_sc_hd__clkbuf_1 _4149_ (.A(_1141_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _4150_ (.A0(net181),
    .A1(\core_0.decode.i_imm_pass[12] ),
    .S(_1133_),
    .X(_1142_));
 sky130_fd_sc_hd__clkbuf_1 _4151_ (.A(_1142_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _4152_ (.A0(net182),
    .A1(\core_0.decode.i_imm_pass[13] ),
    .S(_1133_),
    .X(_1143_));
 sky130_fd_sc_hd__clkbuf_1 _4153_ (.A(_1143_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _4154_ (.A0(net183),
    .A1(\core_0.decode.i_imm_pass[14] ),
    .S(_0913_),
    .X(_1144_));
 sky130_fd_sc_hd__clkbuf_1 _4155_ (.A(_1144_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _4156_ (.A0(net184),
    .A1(\core_0.decode.i_imm_pass[15] ),
    .S(_0913_),
    .X(_1145_));
 sky130_fd_sc_hd__clkbuf_1 _4157_ (.A(_1145_),
    .X(_0054_));
 sky130_fd_sc_hd__clkbuf_4 _4158_ (.A(\core_0.dec_mem_access ),
    .X(_1146_));
 sky130_fd_sc_hd__or2_1 _4159_ (.A(_0976_),
    .B(_1087_),
    .X(_1147_));
 sky130_fd_sc_hd__a22o_1 _4160_ (.A1(_1146_),
    .A2(_1114_),
    .B1(_0952_),
    .B2(_1147_),
    .X(_0055_));
 sky130_fd_sc_hd__a22o_1 _4161_ (.A1(\core_0.dec_mem_we ),
    .A2(_0954_),
    .B1(_0952_),
    .B2(_1107_),
    .X(_0056_));
 sky130_fd_sc_hd__or4_1 _4162_ (.A(_0965_),
    .B(_0979_),
    .C(_1000_),
    .D(_1079_),
    .X(_1148_));
 sky130_fd_sc_hd__or4_2 _4163_ (.A(_0994_),
    .B(_1083_),
    .C(_1100_),
    .D(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__or2_1 _4164_ (.A(\core_0.dec_used_operands[0] ),
    .B(_0909_),
    .X(_1150_));
 sky130_fd_sc_hd__o311a_1 _4165_ (.A1(_1097_),
    .A2(_1111_),
    .A3(_1149_),
    .B1(_1150_),
    .C1(_1075_),
    .X(_0057_));
 sky130_fd_sc_hd__o21ba_1 _4166_ (.A1(_1108_),
    .A2(_1111_),
    .B1_N(_1149_),
    .X(_1151_));
 sky130_fd_sc_hd__a22o_1 _4167_ (.A1(\core_0.dec_used_operands[1] ),
    .A2(_0954_),
    .B1(_1151_),
    .B2(_1075_),
    .X(_0058_));
 sky130_fd_sc_hd__a22o_1 _4168_ (.A1(\core_0.dec_sreg_load ),
    .A2(_0954_),
    .B1(_0952_),
    .B2(_1116_),
    .X(_0059_));
 sky130_fd_sc_hd__clkbuf_8 _4169_ (.A(\core_0.dec_sreg_store ),
    .X(_1152_));
 sky130_fd_sc_hd__a22o_1 _4170_ (.A1(_1152_),
    .A2(_0954_),
    .B1(_0952_),
    .B2(_1106_),
    .X(_0060_));
 sky130_fd_sc_hd__inv_2 _4171_ (.A(_0941_),
    .Y(_1153_));
 sky130_fd_sc_hd__a32o_1 _4172_ (.A1(_0952_),
    .A2(_0935_),
    .A3(_1153_),
    .B1(_0910_),
    .B2(\core_0.dec_sreg_jal_over ),
    .X(_0061_));
 sky130_fd_sc_hd__clkbuf_4 _4173_ (.A(_1038_),
    .X(_1154_));
 sky130_fd_sc_hd__a2bb2o_1 _4174_ (.A1_N(_1128_),
    .A2_N(_1073_),
    .B1(_0911_),
    .B2(_1154_),
    .X(_0062_));
 sky130_fd_sc_hd__nor2_1 _4175_ (.A(_0918_),
    .B(_0939_),
    .Y(_1155_));
 sky130_fd_sc_hd__a22o_1 _4176_ (.A1(\core_0.dec_sys ),
    .A2(_0954_),
    .B1(_0952_),
    .B2(_1155_),
    .X(_0063_));
 sky130_fd_sc_hd__a21o_1 _4177_ (.A1(\core_0.decode.i_instr_l[1] ),
    .A2(_0976_),
    .B1(_1085_),
    .X(_1156_));
 sky130_fd_sc_hd__a22o_1 _4178_ (.A1(\core_0.dec_mem_width ),
    .A2(_0954_),
    .B1(_0952_),
    .B2(_1156_),
    .X(_0064_));
 sky130_fd_sc_hd__a22o_1 _4179_ (.A1(\core_0.dec_mem_long ),
    .A2(_0954_),
    .B1(_0952_),
    .B2(_0976_),
    .X(_0065_));
 sky130_fd_sc_hd__buf_6 _4180_ (.A(_0907_),
    .X(_1157_));
 sky130_fd_sc_hd__or2_2 _4181_ (.A(_1068_),
    .B(_1071_),
    .X(_1158_));
 sky130_fd_sc_hd__nor4_1 _4182_ (.A(_0791_),
    .B(_1157_),
    .C(_1158_),
    .D(_0908_),
    .Y(_0066_));
 sky130_fd_sc_hd__and2_2 _4183_ (.A(net178),
    .B(_1034_),
    .X(_1159_));
 sky130_fd_sc_hd__and3_1 _4184_ (.A(_1032_),
    .B(_1036_),
    .C(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__buf_2 _4185_ (.A(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__clkbuf_4 _4186_ (.A(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__nand2_1 _4187_ (.A(net210),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__nor2_4 _4188_ (.A(_1038_),
    .B(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__nor2_4 _4189_ (.A(_0674_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__buf_4 _4190_ (.A(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__or2_1 _4191_ (.A(_0907_),
    .B(_0674_),
    .X(_1167_));
 sky130_fd_sc_hd__clkbuf_4 _4192_ (.A(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__or2_1 _4193_ (.A(_1154_),
    .B(_1163_),
    .X(_1169_));
 sky130_fd_sc_hd__nor2_1 _4194_ (.A(_0664_),
    .B(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__a211o_1 _4195_ (.A1(\core_0.execute.sreg_priv_control.o_d[0] ),
    .A2(_1166_),
    .B1(_1168_),
    .C1(_1170_),
    .X(_0067_));
 sky130_fd_sc_hd__buf_4 _4196_ (.A(_1164_),
    .X(_1171_));
 sky130_fd_sc_hd__a22o_1 _4197_ (.A1(net201),
    .A2(_1171_),
    .B1(_1166_),
    .B2(\core_0.execute.sreg_data_page ),
    .X(_1172_));
 sky130_fd_sc_hd__and2_1 _4198_ (.A(_1066_),
    .B(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_1 _4199_ (.A(_1173_),
    .X(_0068_));
 sky130_fd_sc_hd__a22o_1 _4200_ (.A1(net203),
    .A2(_1171_),
    .B1(_1166_),
    .B2(\core_0.execute.sreg_long_ptr_en ),
    .X(_1174_));
 sky130_fd_sc_hd__and2_1 _4201_ (.A(_1066_),
    .B(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__clkbuf_1 _4202_ (.A(_1175_),
    .X(_0069_));
 sky130_fd_sc_hd__a22o_1 _4203_ (.A1(net204),
    .A2(_1171_),
    .B1(_1166_),
    .B2(\core_0.execute.sreg_priv_control.o_d[4] ),
    .X(_1176_));
 sky130_fd_sc_hd__and2_1 _4204_ (.A(_1066_),
    .B(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__clkbuf_1 _4205_ (.A(_1177_),
    .X(_0070_));
 sky130_fd_sc_hd__a22o_1 _4206_ (.A1(net205),
    .A2(_1171_),
    .B1(_1166_),
    .B2(\core_0.execute.sreg_priv_control.o_d[5] ),
    .X(_1178_));
 sky130_fd_sc_hd__and2_1 _4207_ (.A(_1066_),
    .B(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__clkbuf_1 _4208_ (.A(_1179_),
    .X(_0071_));
 sky130_fd_sc_hd__a22o_1 _4209_ (.A1(net206),
    .A2(_1171_),
    .B1(_1166_),
    .B2(\core_0.execute.sreg_priv_control.o_d[6] ),
    .X(_1180_));
 sky130_fd_sc_hd__and2_1 _4210_ (.A(_1066_),
    .B(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__clkbuf_1 _4211_ (.A(_1181_),
    .X(_0072_));
 sky130_fd_sc_hd__a22o_1 _4212_ (.A1(net207),
    .A2(_1171_),
    .B1(_1166_),
    .B2(\core_0.execute.sreg_priv_control.o_d[7] ),
    .X(_1182_));
 sky130_fd_sc_hd__and2_1 _4213_ (.A(_1066_),
    .B(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__clkbuf_1 _4214_ (.A(_1183_),
    .X(_0073_));
 sky130_fd_sc_hd__a22o_1 _4215_ (.A1(net208),
    .A2(_1171_),
    .B1(_1166_),
    .B2(\core_0.execute.sreg_priv_control.o_d[8] ),
    .X(_1184_));
 sky130_fd_sc_hd__and2_1 _4216_ (.A(_1066_),
    .B(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__clkbuf_1 _4217_ (.A(_1185_),
    .X(_0074_));
 sky130_fd_sc_hd__a22o_1 _4218_ (.A1(net209),
    .A2(_1171_),
    .B1(_1166_),
    .B2(\core_0.execute.sreg_priv_control.o_d[9] ),
    .X(_1186_));
 sky130_fd_sc_hd__and2_1 _4219_ (.A(_1066_),
    .B(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__clkbuf_1 _4220_ (.A(_1187_),
    .X(_0075_));
 sky130_fd_sc_hd__a22o_1 _4221_ (.A1(net195),
    .A2(_1171_),
    .B1(_1166_),
    .B2(\core_0.execute.sreg_priv_control.o_d[10] ),
    .X(_1188_));
 sky130_fd_sc_hd__and2_1 _4222_ (.A(_1066_),
    .B(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__clkbuf_1 _4223_ (.A(_1189_),
    .X(_0076_));
 sky130_fd_sc_hd__buf_4 _4224_ (.A(_0995_),
    .X(_1190_));
 sky130_fd_sc_hd__a22o_1 _4225_ (.A1(net196),
    .A2(_1171_),
    .B1(_1165_),
    .B2(\core_0.execute.sreg_priv_control.o_d[11] ),
    .X(_1191_));
 sky130_fd_sc_hd__and2_1 _4226_ (.A(_1190_),
    .B(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_1 _4227_ (.A(_1192_),
    .X(_0077_));
 sky130_fd_sc_hd__a22o_1 _4228_ (.A1(net197),
    .A2(_1164_),
    .B1(_1165_),
    .B2(\core_0.execute.sreg_priv_control.o_d[12] ),
    .X(_1193_));
 sky130_fd_sc_hd__and2_1 _4229_ (.A(_1190_),
    .B(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__clkbuf_1 _4230_ (.A(_1194_),
    .X(_0078_));
 sky130_fd_sc_hd__a22o_1 _4231_ (.A1(net198),
    .A2(_1164_),
    .B1(_1165_),
    .B2(\core_0.execute.sreg_priv_control.o_d[13] ),
    .X(_1195_));
 sky130_fd_sc_hd__and2_1 _4232_ (.A(_1190_),
    .B(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__clkbuf_1 _4233_ (.A(_1196_),
    .X(_0079_));
 sky130_fd_sc_hd__a22o_1 _4234_ (.A1(net199),
    .A2(_1164_),
    .B1(_1165_),
    .B2(\core_0.execute.sreg_priv_control.o_d[14] ),
    .X(_1197_));
 sky130_fd_sc_hd__and2_1 _4235_ (.A(_1190_),
    .B(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__clkbuf_1 _4236_ (.A(_1198_),
    .X(_0080_));
 sky130_fd_sc_hd__a22o_1 _4237_ (.A1(net200),
    .A2(_1164_),
    .B1(_1165_),
    .B2(\core_0.execute.sreg_priv_control.o_d[15] ),
    .X(_1199_));
 sky130_fd_sc_hd__and2_1 _4238_ (.A(_1190_),
    .B(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__clkbuf_1 _4239_ (.A(_1200_),
    .X(_0081_));
 sky130_fd_sc_hd__buf_2 _4240_ (.A(\core_0.execute.alu_mul_div.cbit[3] ),
    .X(_1201_));
 sky130_fd_sc_hd__buf_4 _4241_ (.A(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__clkinv_2 _4242_ (.A(\core_0.execute.alu_mul_div.cbit[2] ),
    .Y(_1203_));
 sky130_fd_sc_hd__clkbuf_4 _4243_ (.A(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__buf_4 _4244_ (.A(\core_0.execute.alu_mul_div.cbit[0] ),
    .X(_1205_));
 sky130_fd_sc_hd__clkbuf_4 _4245_ (.A(\core_0.execute.alu_mul_div.cbit[1] ),
    .X(_1206_));
 sky130_fd_sc_hd__buf_4 _4246_ (.A(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__nand2_1 _4247_ (.A(_1205_),
    .B(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__nor2_2 _4248_ (.A(_1204_),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__nand2_4 _4249_ (.A(_1202_),
    .B(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__nor2_1 _4250_ (.A(\core_0.execute.alu_mul_div.comp ),
    .B(_0744_),
    .Y(_1211_));
 sky130_fd_sc_hd__nor4_4 _4251_ (.A(_0791_),
    .B(_0907_),
    .C(_0694_),
    .D(_1211_),
    .Y(_1212_));
 sky130_fd_sc_hd__o21a_1 _4252_ (.A1(_0744_),
    .A2(_1210_),
    .B1(_1212_),
    .X(_0082_));
 sky130_fd_sc_hd__inv_2 _4253_ (.A(_1024_),
    .Y(_1213_));
 sky130_fd_sc_hd__or4b_1 _4254_ (.A(net71),
    .B(_0748_),
    .C(_1213_),
    .D_N(net70),
    .X(_1214_));
 sky130_fd_sc_hd__clkbuf_4 _4255_ (.A(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__buf_4 _4256_ (.A(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__mux2_1 _4257_ (.A0(net38),
    .A1(\core_0.fetch.out_buffer_data_instr[0] ),
    .S(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__clkbuf_1 _4258_ (.A(_1217_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _4259_ (.A0(net49),
    .A1(\core_0.fetch.out_buffer_data_instr[1] ),
    .S(_1216_),
    .X(_1218_));
 sky130_fd_sc_hd__clkbuf_1 _4260_ (.A(_1218_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _4261_ (.A0(net60),
    .A1(\core_0.fetch.out_buffer_data_instr[2] ),
    .S(_1216_),
    .X(_1219_));
 sky130_fd_sc_hd__clkbuf_1 _4262_ (.A(_1219_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(net63),
    .A1(\core_0.fetch.out_buffer_data_instr[3] ),
    .S(_1216_),
    .X(_1220_));
 sky130_fd_sc_hd__clkbuf_1 _4264_ (.A(_1220_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(net64),
    .A1(\core_0.fetch.out_buffer_data_instr[4] ),
    .S(_1216_),
    .X(_1221_));
 sky130_fd_sc_hd__clkbuf_1 _4266_ (.A(_1221_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _4267_ (.A0(net65),
    .A1(\core_0.fetch.out_buffer_data_instr[5] ),
    .S(_1216_),
    .X(_1222_));
 sky130_fd_sc_hd__clkbuf_1 _4268_ (.A(_1222_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _4269_ (.A0(net66),
    .A1(\core_0.fetch.out_buffer_data_instr[6] ),
    .S(_1216_),
    .X(_1223_));
 sky130_fd_sc_hd__clkbuf_1 _4270_ (.A(_1223_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _4271_ (.A0(net67),
    .A1(\core_0.fetch.out_buffer_data_instr[7] ),
    .S(_1216_),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_1 _4272_ (.A(_1224_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _4273_ (.A0(net68),
    .A1(\core_0.fetch.out_buffer_data_instr[8] ),
    .S(_1216_),
    .X(_1225_));
 sky130_fd_sc_hd__clkbuf_1 _4274_ (.A(_1225_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _4275_ (.A0(net69),
    .A1(\core_0.fetch.out_buffer_data_instr[9] ),
    .S(_1216_),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_1 _4276_ (.A(_1226_),
    .X(_0092_));
 sky130_fd_sc_hd__buf_4 _4277_ (.A(_1215_),
    .X(_1227_));
 sky130_fd_sc_hd__mux2_1 _4278_ (.A0(net39),
    .A1(\core_0.fetch.out_buffer_data_instr[10] ),
    .S(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__clkbuf_1 _4279_ (.A(_1228_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _4280_ (.A0(net40),
    .A1(\core_0.fetch.out_buffer_data_instr[11] ),
    .S(_1227_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _4281_ (.A(_1229_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _4282_ (.A0(net41),
    .A1(\core_0.fetch.out_buffer_data_instr[12] ),
    .S(_1227_),
    .X(_1230_));
 sky130_fd_sc_hd__clkbuf_1 _4283_ (.A(_1230_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _4284_ (.A0(net42),
    .A1(\core_0.fetch.out_buffer_data_instr[13] ),
    .S(_1227_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _4285_ (.A(_1231_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _4286_ (.A0(net43),
    .A1(\core_0.fetch.out_buffer_data_instr[14] ),
    .S(_1227_),
    .X(_1232_));
 sky130_fd_sc_hd__clkbuf_1 _4287_ (.A(_1232_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(net44),
    .A1(\core_0.fetch.out_buffer_data_instr[15] ),
    .S(_1227_),
    .X(_1233_));
 sky130_fd_sc_hd__clkbuf_1 _4289_ (.A(_1233_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(net45),
    .A1(\core_0.fetch.out_buffer_data_instr[16] ),
    .S(_1227_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _4291_ (.A(_1234_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(net46),
    .A1(\core_0.fetch.out_buffer_data_instr[17] ),
    .S(_1227_),
    .X(_1235_));
 sky130_fd_sc_hd__clkbuf_1 _4293_ (.A(_1235_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _4294_ (.A0(net47),
    .A1(\core_0.fetch.out_buffer_data_instr[18] ),
    .S(_1227_),
    .X(_1236_));
 sky130_fd_sc_hd__clkbuf_1 _4295_ (.A(_1236_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(net48),
    .A1(\core_0.fetch.out_buffer_data_instr[19] ),
    .S(_1227_),
    .X(_1237_));
 sky130_fd_sc_hd__clkbuf_1 _4297_ (.A(_1237_),
    .X(_0102_));
 sky130_fd_sc_hd__buf_4 _4298_ (.A(_1215_),
    .X(_1238_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(net50),
    .A1(\core_0.fetch.out_buffer_data_instr[20] ),
    .S(_1238_),
    .X(_1239_));
 sky130_fd_sc_hd__clkbuf_1 _4300_ (.A(_1239_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _4301_ (.A0(net51),
    .A1(\core_0.fetch.out_buffer_data_instr[21] ),
    .S(_1238_),
    .X(_1240_));
 sky130_fd_sc_hd__clkbuf_1 _4302_ (.A(_1240_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _4303_ (.A0(net52),
    .A1(\core_0.fetch.out_buffer_data_instr[22] ),
    .S(_1238_),
    .X(_1241_));
 sky130_fd_sc_hd__clkbuf_1 _4304_ (.A(_1241_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _4305_ (.A0(net53),
    .A1(\core_0.fetch.out_buffer_data_instr[23] ),
    .S(_1238_),
    .X(_1242_));
 sky130_fd_sc_hd__clkbuf_1 _4306_ (.A(_1242_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(net54),
    .A1(\core_0.fetch.out_buffer_data_instr[24] ),
    .S(_1238_),
    .X(_1243_));
 sky130_fd_sc_hd__clkbuf_1 _4308_ (.A(_1243_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(net55),
    .A1(\core_0.fetch.out_buffer_data_instr[25] ),
    .S(_1238_),
    .X(_1244_));
 sky130_fd_sc_hd__clkbuf_1 _4310_ (.A(_1244_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(net56),
    .A1(\core_0.fetch.out_buffer_data_instr[26] ),
    .S(_1238_),
    .X(_1245_));
 sky130_fd_sc_hd__clkbuf_1 _4312_ (.A(_1245_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(net57),
    .A1(\core_0.fetch.out_buffer_data_instr[27] ),
    .S(_1238_),
    .X(_1246_));
 sky130_fd_sc_hd__clkbuf_1 _4314_ (.A(_1246_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _4315_ (.A0(net58),
    .A1(\core_0.fetch.out_buffer_data_instr[28] ),
    .S(_1238_),
    .X(_1247_));
 sky130_fd_sc_hd__clkbuf_1 _4316_ (.A(_1247_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _4317_ (.A0(net59),
    .A1(\core_0.fetch.out_buffer_data_instr[29] ),
    .S(_1238_),
    .X(_1248_));
 sky130_fd_sc_hd__clkbuf_1 _4318_ (.A(_1248_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _4319_ (.A0(net61),
    .A1(\core_0.fetch.out_buffer_data_instr[30] ),
    .S(_1215_),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_1 _4320_ (.A(_1249_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(net62),
    .A1(\core_0.fetch.out_buffer_data_instr[31] ),
    .S(_1215_),
    .X(_1250_));
 sky130_fd_sc_hd__clkbuf_1 _4322_ (.A(_1250_),
    .X(_0114_));
 sky130_fd_sc_hd__a21oi_1 _4323_ (.A1(net70),
    .A2(_1024_),
    .B1(_0670_),
    .Y(_1251_));
 sky130_fd_sc_hd__nor4_4 _4324_ (.A(_0791_),
    .B(_1157_),
    .C(_0748_),
    .D(_1251_),
    .Y(_0115_));
 sky130_fd_sc_hd__buf_2 _4325_ (.A(_0788_),
    .X(_1252_));
 sky130_fd_sc_hd__or3_1 _4326_ (.A(_0812_),
    .B(_1122_),
    .C(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__a21bo_1 _4327_ (.A1(net177),
    .A2(net161),
    .B1_N(_1253_),
    .X(_0116_));
 sky130_fd_sc_hd__buf_2 _4328_ (.A(_0907_),
    .X(_1254_));
 sky130_fd_sc_hd__or3_1 _4329_ (.A(_0811_),
    .B(_1254_),
    .C(_1252_),
    .X(_1255_));
 sky130_fd_sc_hd__a21bo_1 _4330_ (.A1(net177),
    .A2(net168),
    .B1_N(_1255_),
    .X(_0117_));
 sky130_fd_sc_hd__or3_1 _4331_ (.A(_0810_),
    .B(_1254_),
    .C(_1252_),
    .X(_1256_));
 sky130_fd_sc_hd__a21bo_1 _4332_ (.A1(net177),
    .A2(net169),
    .B1_N(_1256_),
    .X(_0118_));
 sky130_fd_sc_hd__or3_1 _4333_ (.A(_0809_),
    .B(_1254_),
    .C(_1252_),
    .X(_1257_));
 sky130_fd_sc_hd__a21bo_1 _4334_ (.A1(net177),
    .A2(net170),
    .B1_N(_1257_),
    .X(_0119_));
 sky130_fd_sc_hd__or3_1 _4335_ (.A(_0808_),
    .B(_1254_),
    .C(_1252_),
    .X(_1258_));
 sky130_fd_sc_hd__a21bo_1 _4336_ (.A1(net177),
    .A2(net171),
    .B1_N(_1258_),
    .X(_0120_));
 sky130_fd_sc_hd__or3_1 _4337_ (.A(_0807_),
    .B(_1254_),
    .C(_1252_),
    .X(_1259_));
 sky130_fd_sc_hd__a21bo_1 _4338_ (.A1(net177),
    .A2(net172),
    .B1_N(_1259_),
    .X(_0121_));
 sky130_fd_sc_hd__or3_1 _4339_ (.A(_0805_),
    .B(_1254_),
    .C(_1252_),
    .X(_1260_));
 sky130_fd_sc_hd__a21bo_1 _4340_ (.A1(net177),
    .A2(net173),
    .B1_N(_1260_),
    .X(_0122_));
 sky130_fd_sc_hd__or3_1 _4341_ (.A(_0806_),
    .B(_1254_),
    .C(_1252_),
    .X(_1261_));
 sky130_fd_sc_hd__a21bo_1 _4342_ (.A1(net177),
    .A2(net174),
    .B1_N(_1261_),
    .X(_0123_));
 sky130_fd_sc_hd__or3_1 _4343_ (.A(_0821_),
    .B(_1254_),
    .C(_1252_),
    .X(_1262_));
 sky130_fd_sc_hd__a21bo_1 _4344_ (.A1(_0790_),
    .A2(net175),
    .B1_N(_1262_),
    .X(_0124_));
 sky130_fd_sc_hd__or3b_1 _4345_ (.A(_1122_),
    .B(_0788_),
    .C_N(\core_0.fetch.prev_request_pc[9] ),
    .X(_1263_));
 sky130_fd_sc_hd__a21bo_1 _4346_ (.A1(_0790_),
    .A2(net176),
    .B1_N(_1263_),
    .X(_0125_));
 sky130_fd_sc_hd__or3_1 _4347_ (.A(_0800_),
    .B(_1254_),
    .C(_0788_),
    .X(_1264_));
 sky130_fd_sc_hd__a21bo_1 _4348_ (.A1(_0790_),
    .A2(net162),
    .B1_N(_1264_),
    .X(_0126_));
 sky130_fd_sc_hd__or3b_1 _4349_ (.A(_1122_),
    .B(_0788_),
    .C_N(\core_0.fetch.prev_request_pc[11] ),
    .X(_1265_));
 sky130_fd_sc_hd__a21bo_1 _4350_ (.A1(_0790_),
    .A2(net163),
    .B1_N(_1265_),
    .X(_0127_));
 sky130_fd_sc_hd__or3_1 _4351_ (.A(_0797_),
    .B(_1254_),
    .C(_0788_),
    .X(_1266_));
 sky130_fd_sc_hd__a21bo_1 _4352_ (.A1(_0790_),
    .A2(net164),
    .B1_N(_1266_),
    .X(_0128_));
 sky130_fd_sc_hd__or3_1 _4353_ (.A(_0798_),
    .B(_0907_),
    .C(_0788_),
    .X(_1267_));
 sky130_fd_sc_hd__a21bo_1 _4354_ (.A1(_0790_),
    .A2(net165),
    .B1_N(_1267_),
    .X(_0129_));
 sky130_fd_sc_hd__or3_1 _4355_ (.A(_0794_),
    .B(_0907_),
    .C(_0788_),
    .X(_1268_));
 sky130_fd_sc_hd__a21bo_1 _4356_ (.A1(_0790_),
    .A2(net166),
    .B1_N(_1268_),
    .X(_0130_));
 sky130_fd_sc_hd__or3b_1 _4357_ (.A(_1122_),
    .B(_0788_),
    .C_N(\core_0.fetch.prev_request_pc[15] ),
    .X(_1269_));
 sky130_fd_sc_hd__a21bo_1 _4358_ (.A1(_0790_),
    .A2(net167),
    .B1_N(_1269_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _4359_ (.A0(\core_0.fetch.current_req_branch_pred ),
    .A1(\core_0.fetch.out_buffer_data_pred ),
    .S(_1215_),
    .X(_1270_));
 sky130_fd_sc_hd__clkbuf_1 _4360_ (.A(_1270_),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_4 _4361_ (.A(_1025_),
    .X(_1271_));
 sky130_fd_sc_hd__mux2_1 _4362_ (.A0(_0751_),
    .A1(\core_0.decode.i_instr_l[0] ),
    .S(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__clkbuf_1 _4363_ (.A(_1272_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _4364_ (.A0(_0752_),
    .A1(\core_0.decode.i_instr_l[1] ),
    .S(_1271_),
    .X(_1273_));
 sky130_fd_sc_hd__clkbuf_1 _4365_ (.A(_1273_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _4366_ (.A0(_0754_),
    .A1(\core_0.decode.i_instr_l[2] ),
    .S(_1271_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _4367_ (.A(_1274_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _4368_ (.A0(_0755_),
    .A1(\core_0.decode.i_instr_l[3] ),
    .S(_1271_),
    .X(_1275_));
 sky130_fd_sc_hd__clkbuf_1 _4369_ (.A(_1275_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _4370_ (.A0(_0785_),
    .A1(\core_0.decode.i_instr_l[4] ),
    .S(_1271_),
    .X(_1276_));
 sky130_fd_sc_hd__clkbuf_1 _4371_ (.A(_1276_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _4372_ (.A0(_0750_),
    .A1(\core_0.decode.i_instr_l[5] ),
    .S(_1271_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_1 _4373_ (.A(_1277_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _4374_ (.A0(_0749_),
    .A1(\core_0.decode.i_instr_l[6] ),
    .S(_1271_),
    .X(_1278_));
 sky130_fd_sc_hd__clkbuf_1 _4375_ (.A(_1278_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _4376_ (.A0(_0835_),
    .A1(\core_0.decode.i_instr_l[7] ),
    .S(_1271_),
    .X(_1279_));
 sky130_fd_sc_hd__clkbuf_1 _4377_ (.A(_1279_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _4378_ (.A0(_0837_),
    .A1(\core_0.decode.i_instr_l[8] ),
    .S(_1271_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _4379_ (.A(_1280_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _4380_ (.A0(_0834_),
    .A1(\core_0.decode.i_instr_l[9] ),
    .S(_1271_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_1 _4381_ (.A(_1281_),
    .X(_0142_));
 sky130_fd_sc_hd__buf_4 _4382_ (.A(_1025_),
    .X(_1282_));
 sky130_fd_sc_hd__mux2_1 _4383_ (.A0(_0836_),
    .A1(\core_0.decode.i_instr_l[10] ),
    .S(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__clkbuf_1 _4384_ (.A(_1283_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _4385_ (.A0(net40),
    .A1(\core_0.fetch.out_buffer_data_instr[11] ),
    .S(_0670_),
    .X(_1284_));
 sky130_fd_sc_hd__mux2_1 _4386_ (.A0(_1284_),
    .A1(\core_0.decode.i_instr_l[11] ),
    .S(_1282_),
    .X(_1285_));
 sky130_fd_sc_hd__clkbuf_1 _4387_ (.A(_1285_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _4388_ (.A0(net41),
    .A1(\core_0.fetch.out_buffer_data_instr[12] ),
    .S(_0670_),
    .X(_1286_));
 sky130_fd_sc_hd__mux2_1 _4389_ (.A0(_1286_),
    .A1(\core_0.decode.i_instr_l[12] ),
    .S(_1282_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_1 _4390_ (.A(_1287_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _4391_ (.A0(net42),
    .A1(\core_0.fetch.out_buffer_data_instr[13] ),
    .S(_0670_),
    .X(_1288_));
 sky130_fd_sc_hd__mux2_1 _4392_ (.A0(_1288_),
    .A1(\core_0.decode.i_instr_l[13] ),
    .S(_1282_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _4393_ (.A(_1289_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _4394_ (.A0(net43),
    .A1(\core_0.fetch.out_buffer_data_instr[14] ),
    .S(_0670_),
    .X(_1290_));
 sky130_fd_sc_hd__mux2_1 _4395_ (.A0(_1290_),
    .A1(\core_0.decode.i_instr_l[14] ),
    .S(_1282_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _4396_ (.A(_1291_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _4397_ (.A0(net44),
    .A1(\core_0.fetch.out_buffer_data_instr[15] ),
    .S(_0670_),
    .X(_1292_));
 sky130_fd_sc_hd__mux2_1 _4398_ (.A0(_1292_),
    .A1(\core_0.decode.i_instr_l[15] ),
    .S(_1282_),
    .X(_1293_));
 sky130_fd_sc_hd__clkbuf_1 _4399_ (.A(_1293_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _4400_ (.A0(_0771_),
    .A1(\core_0.decode.i_imm_pass[0] ),
    .S(_1282_),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _4401_ (.A(_1294_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _4402_ (.A0(_0759_),
    .A1(\core_0.decode.i_imm_pass[1] ),
    .S(_1282_),
    .X(_1295_));
 sky130_fd_sc_hd__clkbuf_1 _4403_ (.A(_1295_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _4404_ (.A0(_0766_),
    .A1(\core_0.decode.i_imm_pass[2] ),
    .S(_1282_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _4405_ (.A(_1296_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _4406_ (.A0(_0761_),
    .A1(\core_0.decode.i_imm_pass[3] ),
    .S(_1282_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_1 _4407_ (.A(_1297_),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_4 _4408_ (.A(_1025_),
    .X(_1298_));
 sky130_fd_sc_hd__mux2_1 _4409_ (.A0(_0763_),
    .A1(\core_0.decode.i_imm_pass[4] ),
    .S(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__clkbuf_1 _4410_ (.A(_1299_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _4411_ (.A0(_0772_),
    .A1(\core_0.decode.i_imm_pass[5] ),
    .S(_1298_),
    .X(_1300_));
 sky130_fd_sc_hd__clkbuf_1 _4412_ (.A(_1300_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _4413_ (.A0(_0774_),
    .A1(\core_0.decode.i_imm_pass[6] ),
    .S(_1298_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_1 _4414_ (.A(_1301_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _4415_ (.A0(_0765_),
    .A1(\core_0.decode.i_imm_pass[7] ),
    .S(_1298_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _4416_ (.A(_1302_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _4417_ (.A0(_0758_),
    .A1(\core_0.decode.i_imm_pass[8] ),
    .S(_1298_),
    .X(_1303_));
 sky130_fd_sc_hd__clkbuf_1 _4418_ (.A(_1303_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _4419_ (.A0(_0778_),
    .A1(\core_0.decode.i_imm_pass[9] ),
    .S(_1298_),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_1 _4420_ (.A(_1304_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _4421_ (.A0(_0760_),
    .A1(\core_0.decode.i_imm_pass[10] ),
    .S(_1298_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_1 _4422_ (.A(_1305_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _4423_ (.A0(_0776_),
    .A1(\core_0.decode.i_imm_pass[11] ),
    .S(_1298_),
    .X(_1306_));
 sky130_fd_sc_hd__clkbuf_1 _4424_ (.A(_1306_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _4425_ (.A0(_0768_),
    .A1(\core_0.decode.i_imm_pass[12] ),
    .S(_1298_),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_1 _4426_ (.A(_1307_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _4427_ (.A0(_0779_),
    .A1(\core_0.decode.i_imm_pass[13] ),
    .S(_1298_),
    .X(_1308_));
 sky130_fd_sc_hd__clkbuf_1 _4428_ (.A(_1308_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _4429_ (.A0(_0764_),
    .A1(\core_0.decode.i_imm_pass[14] ),
    .S(_1025_),
    .X(_1309_));
 sky130_fd_sc_hd__clkbuf_1 _4430_ (.A(_1309_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _4431_ (.A0(_0770_),
    .A1(\core_0.decode.i_imm_pass[15] ),
    .S(_1025_),
    .X(_1310_));
 sky130_fd_sc_hd__clkbuf_1 _4432_ (.A(_1310_),
    .X(_0164_));
 sky130_fd_sc_hd__nor2_1 _4433_ (.A(_1122_),
    .B(net70),
    .Y(_1311_));
 sky130_fd_sc_hd__a21o_1 _4434_ (.A1(\core_0.fetch.dbg_out ),
    .A2(_1311_),
    .B1(net177),
    .X(_0165_));
 sky130_fd_sc_hd__o211a_1 _4435_ (.A1(\core_0.fetch.flush_event_invalidate ),
    .A2(\core_0.fetch.dbg_out ),
    .B1(_1213_),
    .C1(_1311_),
    .X(_0166_));
 sky130_fd_sc_hd__and3b_1 _4436_ (.A_N(_1252_),
    .B(_0862_),
    .C(_0995_),
    .X(_1312_));
 sky130_fd_sc_hd__clkbuf_1 _4437_ (.A(_1312_),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_1 _4438_ (.A(_1122_),
    .X(_1313_));
 sky130_fd_sc_hd__clkbuf_1 _4439_ (.A(_1313_),
    .X(_0168_));
 sky130_fd_sc_hd__buf_6 _4440_ (.A(_0995_),
    .X(_1314_));
 sky130_fd_sc_hd__buf_4 _4441_ (.A(net37),
    .X(_1315_));
 sky130_fd_sc_hd__clkinv_2 _4442_ (.A(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__clkbuf_4 _4443_ (.A(\core_0.ew_mem_access ),
    .X(_1317_));
 sky130_fd_sc_hd__buf_4 _4444_ (.A(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__mux2_1 _4445_ (.A0(_1316_),
    .A1(_1318_),
    .S(\core_0.ew_submit ),
    .X(_1319_));
 sky130_fd_sc_hd__and3_1 _4446_ (.A(_1314_),
    .B(_0740_),
    .C(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__clkbuf_1 _4447_ (.A(_1320_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _4448_ (.A0(\core_0.fetch.current_req_branch_pred ),
    .A1(\core_0.fetch.out_buffer_data_pred ),
    .S(_0670_),
    .X(_1321_));
 sky130_fd_sc_hd__mux2_1 _4449_ (.A0(\core_0.decode.i_jmp_pred_pass ),
    .A1(_1321_),
    .S(\core_0.fetch.submitable ),
    .X(_1322_));
 sky130_fd_sc_hd__clkbuf_1 _4450_ (.A(_1322_),
    .X(_0170_));
 sky130_fd_sc_hd__and2_1 _4451_ (.A(_1076_),
    .B(net184),
    .X(_1323_));
 sky130_fd_sc_hd__inv_2 _4452_ (.A(\core_0.dec_r_bus_imm ),
    .Y(_1324_));
 sky130_fd_sc_hd__o221a_2 _4453_ (.A1(net94),
    .A2(_0520_),
    .B1(_0529_),
    .B2(_0540_),
    .C1(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__nor2_4 _4454_ (.A(_1323_),
    .B(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__or2_1 _4455_ (.A(\core_0.execute.alu_mul_div.div_cur[15] ),
    .B(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__and2_1 _4456_ (.A(_1076_),
    .B(net183),
    .X(_1328_));
 sky130_fd_sc_hd__buf_6 _4457_ (.A(_1324_),
    .X(_1329_));
 sky130_fd_sc_hd__o311a_2 _4458_ (.A1(_0544_),
    .A2(_0548_),
    .A3(_0551_),
    .B1(_0552_),
    .C1(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__or2_4 _4459_ (.A(_1328_),
    .B(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__clkinv_2 _4460_ (.A(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__o221a_2 _4461_ (.A1(net92),
    .A2(_0521_),
    .B1(_0562_),
    .B2(_0567_),
    .C1(_1329_),
    .X(_1333_));
 sky130_fd_sc_hd__a21oi_4 _4462_ (.A1(_1077_),
    .A2(net182),
    .B1(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__and2_1 _4463_ (.A(\core_0.execute.alu_mul_div.div_cur[13] ),
    .B(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__and2_1 _4464_ (.A(_1076_),
    .B(net181),
    .X(_1336_));
 sky130_fd_sc_hd__o221a_2 _4465_ (.A1(net91),
    .A2(_0521_),
    .B1(_0575_),
    .B2(_0578_),
    .C1(_1329_),
    .X(_1337_));
 sky130_fd_sc_hd__nor2_4 _4466_ (.A(_1336_),
    .B(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__inv_2 _4467_ (.A(net180),
    .Y(_1339_));
 sky130_fd_sc_hd__clkinv_2 _4468_ (.A(net196),
    .Y(_1340_));
 sky130_fd_sc_hd__buf_6 _4469_ (.A(_1329_),
    .X(_1341_));
 sky130_fd_sc_hd__mux2_4 _4470_ (.A0(_1339_),
    .A1(_1340_),
    .S(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__nand2_1 _4471_ (.A(\core_0.execute.alu_mul_div.div_cur[11] ),
    .B(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__mux2_4 _4472_ (.A0(net179),
    .A1(net195),
    .S(_1329_),
    .X(_1344_));
 sky130_fd_sc_hd__clkinv_2 _4473_ (.A(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__and2_1 _4474_ (.A(\core_0.execute.alu_mul_div.div_cur[10] ),
    .B(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__nor2_1 _4475_ (.A(\core_0.execute.alu_mul_div.div_cur[10] ),
    .B(_1345_),
    .Y(_1347_));
 sky130_fd_sc_hd__nor2_1 _4476_ (.A(_1346_),
    .B(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__inv_2 _4477_ (.A(net193),
    .Y(_1349_));
 sky130_fd_sc_hd__mux2_4 _4478_ (.A0(_1349_),
    .A1(_0598_),
    .S(_1341_),
    .X(_1350_));
 sky130_fd_sc_hd__or2_1 _4479_ (.A(\core_0.execute.alu_mul_div.div_cur[9] ),
    .B(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__o211a_2 _4480_ (.A1(_0608_),
    .A2(_0611_),
    .B1(_0612_),
    .C1(_1329_),
    .X(_1352_));
 sky130_fd_sc_hd__a21oi_4 _4481_ (.A1(_1077_),
    .A2(net191),
    .B1(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__or2_1 _4482_ (.A(\core_0.execute.alu_mul_div.div_cur[7] ),
    .B(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__and2_1 _4483_ (.A(_1076_),
    .B(net190),
    .X(_1355_));
 sky130_fd_sc_hd__o311a_1 _4484_ (.A1(_0617_),
    .A2(_0618_),
    .A3(_0619_),
    .B1(_0620_),
    .C1(_1329_),
    .X(_1356_));
 sky130_fd_sc_hd__or2_4 _4485_ (.A(_1355_),
    .B(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__and2b_1 _4486_ (.A_N(_1357_),
    .B(\core_0.execute.alu_mul_div.div_cur[6] ),
    .X(_1358_));
 sky130_fd_sc_hd__and2b_1 _4487_ (.A_N(\core_0.execute.alu_mul_div.div_cur[6] ),
    .B(_1357_),
    .X(_1359_));
 sky130_fd_sc_hd__nor2_1 _4488_ (.A(_1358_),
    .B(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__nor2_2 _4489_ (.A(_1341_),
    .B(net189),
    .Y(_1361_));
 sky130_fd_sc_hd__a21o_4 _4490_ (.A1(_1341_),
    .A2(_0627_),
    .B1(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__or2_1 _4491_ (.A(\core_0.execute.alu_mul_div.div_cur[5] ),
    .B(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__nand2_1 _4492_ (.A(_1076_),
    .B(net188),
    .Y(_1364_));
 sky130_fd_sc_hd__o21a_4 _4493_ (.A1(_1077_),
    .A2(_0633_),
    .B1(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__and2_1 _4494_ (.A(\core_0.execute.alu_mul_div.div_cur[4] ),
    .B(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__nor2_1 _4495_ (.A(\core_0.execute.alu_mul_div.div_cur[4] ),
    .B(_1365_),
    .Y(_1367_));
 sky130_fd_sc_hd__nor2_1 _4496_ (.A(_1366_),
    .B(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__inv_2 _4497_ (.A(net187),
    .Y(_1369_));
 sky130_fd_sc_hd__mux2_4 _4498_ (.A0(_1369_),
    .A1(_0639_),
    .S(_1341_),
    .X(_1370_));
 sky130_fd_sc_hd__buf_6 _4499_ (.A(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__or2_1 _4500_ (.A(\core_0.execute.alu_mul_div.div_cur[3] ),
    .B(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__or2_1 _4501_ (.A(_1329_),
    .B(net186),
    .X(_1373_));
 sky130_fd_sc_hd__o21ai_4 _4502_ (.A1(_1077_),
    .A2(net202),
    .B1(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__nor2_1 _4503_ (.A(\core_0.execute.alu_mul_div.div_cur[2] ),
    .B(_1374_),
    .Y(_1375_));
 sky130_fd_sc_hd__nand2_8 _4504_ (.A(\core_0.dec_r_bus_imm ),
    .B(net178),
    .Y(_1376_));
 sky130_fd_sc_hd__a211o_4 _4505_ (.A1(_0659_),
    .A2(_0662_),
    .B1(_1076_),
    .C1(_0663_),
    .X(_1377_));
 sky130_fd_sc_hd__a21o_1 _4506_ (.A1(_1376_),
    .A2(_1377_),
    .B1(\core_0.execute.alu_mul_div.div_cur[0] ),
    .X(_1378_));
 sky130_fd_sc_hd__nand2_4 _4507_ (.A(_1076_),
    .B(net185),
    .Y(_1379_));
 sky130_fd_sc_hd__o221ai_4 _4508_ (.A1(net95),
    .A2(_0521_),
    .B1(_0651_),
    .B2(_0654_),
    .C1(_1329_),
    .Y(_1380_));
 sky130_fd_sc_hd__a21o_1 _4509_ (.A1(_1379_),
    .A2(_1380_),
    .B1(\core_0.execute.alu_mul_div.div_cur[1] ),
    .X(_1381_));
 sky130_fd_sc_hd__and3_1 _4510_ (.A(\core_0.execute.alu_mul_div.div_cur[1] ),
    .B(_1379_),
    .C(_1380_),
    .X(_1382_));
 sky130_fd_sc_hd__a21oi_2 _4511_ (.A1(_1378_),
    .A2(_1381_),
    .B1(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__nand2_1 _4512_ (.A(\core_0.execute.alu_mul_div.div_cur[3] ),
    .B(_1370_),
    .Y(_1384_));
 sky130_fd_sc_hd__nand2_1 _4513_ (.A(\core_0.execute.alu_mul_div.div_cur[2] ),
    .B(_1374_),
    .Y(_1385_));
 sky130_fd_sc_hd__o211ai_2 _4514_ (.A1(_1375_),
    .A2(_1383_),
    .B1(_1384_),
    .C1(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__and2_1 _4515_ (.A(\core_0.execute.alu_mul_div.div_cur[5] ),
    .B(_1362_),
    .X(_1387_));
 sky130_fd_sc_hd__a311o_1 _4516_ (.A1(_1368_),
    .A2(_1372_),
    .A3(_1386_),
    .B1(_1366_),
    .C1(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__and2_1 _4517_ (.A(\core_0.execute.alu_mul_div.div_cur[7] ),
    .B(_1353_),
    .X(_1389_));
 sky130_fd_sc_hd__a311o_1 _4518_ (.A1(_1360_),
    .A2(_1363_),
    .A3(_1388_),
    .B1(_1358_),
    .C1(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__mux2_4 _4519_ (.A0(net192),
    .A1(net208),
    .S(_1341_),
    .X(_1391_));
 sky130_fd_sc_hd__inv_2 _4520_ (.A(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__and2_1 _4521_ (.A(\core_0.execute.alu_mul_div.div_cur[8] ),
    .B(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__nor2_1 _4522_ (.A(\core_0.execute.alu_mul_div.div_cur[8] ),
    .B(_1392_),
    .Y(_1394_));
 sky130_fd_sc_hd__nor2_1 _4523_ (.A(_1393_),
    .B(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__and2_1 _4524_ (.A(\core_0.execute.alu_mul_div.div_cur[9] ),
    .B(_1350_),
    .X(_1396_));
 sky130_fd_sc_hd__a311o_1 _4525_ (.A1(_1354_),
    .A2(_1390_),
    .A3(_1395_),
    .B1(_1393_),
    .C1(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__a31o_1 _4526_ (.A1(_1348_),
    .A2(_1351_),
    .A3(_1397_),
    .B1(_1346_),
    .X(_1398_));
 sky130_fd_sc_hd__o21ai_1 _4527_ (.A1(\core_0.execute.alu_mul_div.div_cur[11] ),
    .A2(_1342_),
    .B1(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__or2_2 _4528_ (.A(_1336_),
    .B(_1337_),
    .X(_1400_));
 sky130_fd_sc_hd__xnor2_1 _4529_ (.A(\core_0.execute.alu_mul_div.div_cur[12] ),
    .B(_1400_),
    .Y(_1401_));
 sky130_fd_sc_hd__a21boi_1 _4530_ (.A1(_1343_),
    .A2(_1399_),
    .B1_N(_1401_),
    .Y(_1402_));
 sky130_fd_sc_hd__a21o_1 _4531_ (.A1(\core_0.execute.alu_mul_div.div_cur[12] ),
    .A2(_1338_),
    .B1(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__xnor2_1 _4532_ (.A(\core_0.execute.alu_mul_div.div_cur[14] ),
    .B(_1331_),
    .Y(_1404_));
 sky130_fd_sc_hd__or2_1 _4533_ (.A(\core_0.execute.alu_mul_div.div_cur[13] ),
    .B(_1334_),
    .X(_1405_));
 sky130_fd_sc_hd__o211a_1 _4534_ (.A1(_1335_),
    .A2(_1403_),
    .B1(_1404_),
    .C1(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__a21o_1 _4535_ (.A1(\core_0.execute.alu_mul_div.div_cur[14] ),
    .A2(_1332_),
    .B1(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__and2_1 _4536_ (.A(\core_0.execute.alu_mul_div.div_cur[15] ),
    .B(_1326_),
    .X(_1408_));
 sky130_fd_sc_hd__a21o_4 _4537_ (.A1(_1327_),
    .A2(_1407_),
    .B1(_1408_),
    .X(_1409_));
 sky130_fd_sc_hd__buf_4 _4538_ (.A(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__buf_2 _4539_ (.A(_0741_),
    .X(_1411_));
 sky130_fd_sc_hd__and2_2 _4540_ (.A(\core_0.execute.alu_mul_div.comp ),
    .B(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__o21a_2 _4541_ (.A1(_1210_),
    .A2(_1410_),
    .B1(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_4 _4542_ (.A(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__o21ai_4 _4543_ (.A1(_1210_),
    .A2(_1409_),
    .B1(_1412_),
    .Y(_1415_));
 sky130_fd_sc_hd__clkbuf_4 _4544_ (.A(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__and2b_1 _4545_ (.A_N(_1382_),
    .B(_1381_),
    .X(_1417_));
 sky130_fd_sc_hd__xor2_1 _4546_ (.A(_1378_),
    .B(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__inv_2 _4547_ (.A(_1376_),
    .Y(_1419_));
 sky130_fd_sc_hd__a211oi_4 _4548_ (.A1(_0659_),
    .A2(_0662_),
    .B1(_1076_),
    .C1(_0663_),
    .Y(_1420_));
 sky130_fd_sc_hd__nor2_4 _4549_ (.A(_1419_),
    .B(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__buf_4 _4550_ (.A(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_4 _4551_ (.A(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__nand2_1 _4552_ (.A(\core_0.execute.alu_mul_div.div_cur[0] ),
    .B(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__and2_1 _4553_ (.A(_1378_),
    .B(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__nand2_1 _4554_ (.A(_1210_),
    .B(_1425_),
    .Y(_1426_));
 sky130_fd_sc_hd__o21a_1 _4555_ (.A1(_1210_),
    .A2(_1418_),
    .B1(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__mux2_1 _4556_ (.A0(\core_0.execute.alu_mul_div.div_cur[0] ),
    .A1(_1427_),
    .S(_1410_),
    .X(_1428_));
 sky130_fd_sc_hd__or2_1 _4557_ (.A(_1416_),
    .B(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__clkbuf_4 _4558_ (.A(_0742_),
    .X(_1430_));
 sky130_fd_sc_hd__o211a_1 _4559_ (.A1(\core_0.execute.alu_mul_div.div_cur[1] ),
    .A2(_1414_),
    .B1(_1429_),
    .C1(_1430_),
    .X(_0171_));
 sky130_fd_sc_hd__buf_4 _4560_ (.A(_1374_),
    .X(_1431_));
 sky130_fd_sc_hd__and2_1 _4561_ (.A(\core_0.execute.alu_mul_div.div_cur[2] ),
    .B(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__nor2_1 _4562_ (.A(_1432_),
    .B(_1375_),
    .Y(_1433_));
 sky130_fd_sc_hd__xnor2_1 _4563_ (.A(_1433_),
    .B(_1383_),
    .Y(_1434_));
 sky130_fd_sc_hd__clkbuf_4 _4564_ (.A(\core_0.execute.alu_mul_div.cbit[2] ),
    .X(_1435_));
 sky130_fd_sc_hd__buf_4 _4565_ (.A(_1435_),
    .X(_1436_));
 sky130_fd_sc_hd__and2_2 _4566_ (.A(_1205_),
    .B(_1207_),
    .X(_1437_));
 sky130_fd_sc_hd__and3_2 _4567_ (.A(_1202_),
    .B(_1436_),
    .C(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__clkbuf_4 _4568_ (.A(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__mux2_1 _4569_ (.A0(_1418_),
    .A1(_1434_),
    .S(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__mux2_1 _4570_ (.A0(\core_0.execute.alu_mul_div.div_cur[1] ),
    .A1(_1440_),
    .S(_1410_),
    .X(_1441_));
 sky130_fd_sc_hd__or2_1 _4571_ (.A(_1416_),
    .B(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__o211a_1 _4572_ (.A1(\core_0.execute.alu_mul_div.div_cur[2] ),
    .A2(_1414_),
    .B1(_1442_),
    .C1(_1430_),
    .X(_0172_));
 sky130_fd_sc_hd__o21ai_1 _4573_ (.A1(_1375_),
    .A2(_1383_),
    .B1(_1385_),
    .Y(_1443_));
 sky130_fd_sc_hd__nand2_1 _4574_ (.A(_1372_),
    .B(_1384_),
    .Y(_1444_));
 sky130_fd_sc_hd__xnor2_1 _4575_ (.A(_1443_),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__mux2_1 _4576_ (.A0(_1434_),
    .A1(_1445_),
    .S(_1439_),
    .X(_1446_));
 sky130_fd_sc_hd__mux2_1 _4577_ (.A0(\core_0.execute.alu_mul_div.div_cur[2] ),
    .A1(_1446_),
    .S(_1410_),
    .X(_1447_));
 sky130_fd_sc_hd__or2_1 _4578_ (.A(_1416_),
    .B(_1447_),
    .X(_1448_));
 sky130_fd_sc_hd__o211a_1 _4579_ (.A1(\core_0.execute.alu_mul_div.div_cur[3] ),
    .A2(_1414_),
    .B1(_1448_),
    .C1(_1430_),
    .X(_0173_));
 sky130_fd_sc_hd__and3_1 _4580_ (.A(_1368_),
    .B(_1372_),
    .C(_1386_),
    .X(_1449_));
 sky130_fd_sc_hd__a21oi_1 _4581_ (.A1(_1372_),
    .A2(_1386_),
    .B1(_1368_),
    .Y(_1450_));
 sky130_fd_sc_hd__nor2_1 _4582_ (.A(_1449_),
    .B(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__mux2_1 _4583_ (.A0(_1445_),
    .A1(_1451_),
    .S(_1439_),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_1 _4584_ (.A0(\core_0.execute.alu_mul_div.div_cur[3] ),
    .A1(_1452_),
    .S(_1410_),
    .X(_1453_));
 sky130_fd_sc_hd__or2_1 _4585_ (.A(_1416_),
    .B(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__o211a_1 _4586_ (.A1(\core_0.execute.alu_mul_div.div_cur[4] ),
    .A2(_1414_),
    .B1(_1454_),
    .C1(_1430_),
    .X(_0174_));
 sky130_fd_sc_hd__or2_1 _4587_ (.A(_1366_),
    .B(_1449_),
    .X(_1455_));
 sky130_fd_sc_hd__and2b_1 _4588_ (.A_N(_1387_),
    .B(_1363_),
    .X(_1456_));
 sky130_fd_sc_hd__xor2_1 _4589_ (.A(_1455_),
    .B(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__mux2_1 _4590_ (.A0(_1451_),
    .A1(_1457_),
    .S(_1439_),
    .X(_1458_));
 sky130_fd_sc_hd__mux2_1 _4591_ (.A0(\core_0.execute.alu_mul_div.div_cur[4] ),
    .A1(_1458_),
    .S(_1410_),
    .X(_1459_));
 sky130_fd_sc_hd__or2_1 _4592_ (.A(_1416_),
    .B(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__o211a_1 _4593_ (.A1(\core_0.execute.alu_mul_div.div_cur[5] ),
    .A2(_1414_),
    .B1(_1460_),
    .C1(_1430_),
    .X(_0175_));
 sky130_fd_sc_hd__and3_1 _4594_ (.A(_1360_),
    .B(_1363_),
    .C(_1388_),
    .X(_1461_));
 sky130_fd_sc_hd__a21oi_1 _4595_ (.A1(_1363_),
    .A2(_1388_),
    .B1(_1360_),
    .Y(_1462_));
 sky130_fd_sc_hd__nor2_1 _4596_ (.A(_1461_),
    .B(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__mux2_1 _4597_ (.A0(_1457_),
    .A1(_1463_),
    .S(_1439_),
    .X(_1464_));
 sky130_fd_sc_hd__mux2_1 _4598_ (.A0(\core_0.execute.alu_mul_div.div_cur[5] ),
    .A1(_1464_),
    .S(_1410_),
    .X(_1465_));
 sky130_fd_sc_hd__or2_1 _4599_ (.A(_1416_),
    .B(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__o211a_1 _4600_ (.A1(\core_0.execute.alu_mul_div.div_cur[6] ),
    .A2(_1414_),
    .B1(_1466_),
    .C1(_1430_),
    .X(_0176_));
 sky130_fd_sc_hd__or2_1 _4601_ (.A(_1358_),
    .B(_1461_),
    .X(_1467_));
 sky130_fd_sc_hd__inv_2 _4602_ (.A(_1354_),
    .Y(_1468_));
 sky130_fd_sc_hd__nor2_1 _4603_ (.A(_1468_),
    .B(_1389_),
    .Y(_1469_));
 sky130_fd_sc_hd__xor2_1 _4604_ (.A(_1467_),
    .B(_1469_),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_1 _4605_ (.A0(_1463_),
    .A1(_1470_),
    .S(_1439_),
    .X(_1471_));
 sky130_fd_sc_hd__mux2_1 _4606_ (.A0(\core_0.execute.alu_mul_div.div_cur[6] ),
    .A1(_1471_),
    .S(_1410_),
    .X(_1472_));
 sky130_fd_sc_hd__or2_1 _4607_ (.A(_1416_),
    .B(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__clkbuf_4 _4608_ (.A(_0742_),
    .X(_1474_));
 sky130_fd_sc_hd__o211a_1 _4609_ (.A1(\core_0.execute.alu_mul_div.div_cur[7] ),
    .A2(_1414_),
    .B1(_1473_),
    .C1(_1474_),
    .X(_0177_));
 sky130_fd_sc_hd__and3_1 _4610_ (.A(_1354_),
    .B(_1390_),
    .C(_1395_),
    .X(_1475_));
 sky130_fd_sc_hd__a21oi_1 _4611_ (.A1(_1354_),
    .A2(_1390_),
    .B1(_1395_),
    .Y(_1476_));
 sky130_fd_sc_hd__nor2_1 _4612_ (.A(_1475_),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__mux2_1 _4613_ (.A0(_1470_),
    .A1(_1477_),
    .S(_1439_),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_1 _4614_ (.A0(\core_0.execute.alu_mul_div.div_cur[7] ),
    .A1(_1478_),
    .S(_1410_),
    .X(_1479_));
 sky130_fd_sc_hd__or2_1 _4615_ (.A(_1416_),
    .B(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__o211a_1 _4616_ (.A1(\core_0.execute.alu_mul_div.div_cur[8] ),
    .A2(_1414_),
    .B1(_1480_),
    .C1(_1474_),
    .X(_0178_));
 sky130_fd_sc_hd__nor2_1 _4617_ (.A(_1393_),
    .B(_1475_),
    .Y(_1481_));
 sky130_fd_sc_hd__mux2_8 _4618_ (.A0(net193),
    .A1(net209),
    .S(_1341_),
    .X(_1482_));
 sky130_fd_sc_hd__xnor2_1 _4619_ (.A(\core_0.execute.alu_mul_div.div_cur[9] ),
    .B(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__xnor2_1 _4620_ (.A(_1481_),
    .B(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__mux2_1 _4621_ (.A0(_1477_),
    .A1(_1484_),
    .S(_1439_),
    .X(_1485_));
 sky130_fd_sc_hd__mux2_1 _4622_ (.A0(\core_0.execute.alu_mul_div.div_cur[8] ),
    .A1(_1485_),
    .S(_1409_),
    .X(_1486_));
 sky130_fd_sc_hd__or2_1 _4623_ (.A(_1416_),
    .B(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__o211a_1 _4624_ (.A1(\core_0.execute.alu_mul_div.div_cur[9] ),
    .A2(_1414_),
    .B1(_1487_),
    .C1(_1474_),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_1 _4625_ (.A(_1351_),
    .B(_1397_),
    .Y(_1488_));
 sky130_fd_sc_hd__xnor2_1 _4626_ (.A(_1348_),
    .B(_1488_),
    .Y(_1489_));
 sky130_fd_sc_hd__mux2_1 _4627_ (.A0(_1484_),
    .A1(_1489_),
    .S(_1439_),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _4628_ (.A0(\core_0.execute.alu_mul_div.div_cur[9] ),
    .A1(_1490_),
    .S(_1409_),
    .X(_1491_));
 sky130_fd_sc_hd__or2_1 _4629_ (.A(_1415_),
    .B(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__o211a_1 _4630_ (.A1(\core_0.execute.alu_mul_div.div_cur[10] ),
    .A2(_1414_),
    .B1(_1492_),
    .C1(_1474_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_8 _4631_ (.A0(net180),
    .A1(net196),
    .S(_1329_),
    .X(_1493_));
 sky130_fd_sc_hd__xor2_2 _4632_ (.A(\core_0.execute.alu_mul_div.div_cur[11] ),
    .B(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__xnor2_1 _4633_ (.A(_1398_),
    .B(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__mux2_1 _4634_ (.A0(_1489_),
    .A1(_1495_),
    .S(_1438_),
    .X(_1496_));
 sky130_fd_sc_hd__mux2_1 _4635_ (.A0(\core_0.execute.alu_mul_div.div_cur[10] ),
    .A1(_1496_),
    .S(_1409_),
    .X(_1497_));
 sky130_fd_sc_hd__or2_1 _4636_ (.A(_1415_),
    .B(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__o211a_1 _4637_ (.A1(\core_0.execute.alu_mul_div.div_cur[11] ),
    .A2(_1413_),
    .B1(_1498_),
    .C1(_1474_),
    .X(_0181_));
 sky130_fd_sc_hd__and3b_1 _4638_ (.A_N(_1401_),
    .B(_1343_),
    .C(_1399_),
    .X(_1499_));
 sky130_fd_sc_hd__nor2_1 _4639_ (.A(_1402_),
    .B(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__mux2_1 _4640_ (.A0(_1495_),
    .A1(_1500_),
    .S(_1438_),
    .X(_1501_));
 sky130_fd_sc_hd__mux2_1 _4641_ (.A0(\core_0.execute.alu_mul_div.div_cur[11] ),
    .A1(_1501_),
    .S(_1409_),
    .X(_1502_));
 sky130_fd_sc_hd__or2_1 _4642_ (.A(_1415_),
    .B(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__o211a_1 _4643_ (.A1(\core_0.execute.alu_mul_div.div_cur[12] ),
    .A2(_1413_),
    .B1(_1503_),
    .C1(_1474_),
    .X(_0182_));
 sky130_fd_sc_hd__inv_2 _4644_ (.A(_1335_),
    .Y(_1504_));
 sky130_fd_sc_hd__nand2_1 _4645_ (.A(_1405_),
    .B(_1504_),
    .Y(_1505_));
 sky130_fd_sc_hd__xnor2_1 _4646_ (.A(_1403_),
    .B(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__mux2_1 _4647_ (.A0(_1500_),
    .A1(_1506_),
    .S(_1438_),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _4648_ (.A0(\core_0.execute.alu_mul_div.div_cur[12] ),
    .A1(_1507_),
    .S(_1409_),
    .X(_1508_));
 sky130_fd_sc_hd__or2_1 _4649_ (.A(_1415_),
    .B(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__o211a_1 _4650_ (.A1(\core_0.execute.alu_mul_div.div_cur[13] ),
    .A2(_1413_),
    .B1(_1509_),
    .C1(_1474_),
    .X(_0183_));
 sky130_fd_sc_hd__o21a_1 _4651_ (.A1(_1335_),
    .A2(_1403_),
    .B1(_1405_),
    .X(_1510_));
 sky130_fd_sc_hd__nor2_1 _4652_ (.A(_1404_),
    .B(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__nor2_1 _4653_ (.A(_1406_),
    .B(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__mux2_1 _4654_ (.A0(_1506_),
    .A1(_1512_),
    .S(_1438_),
    .X(_1513_));
 sky130_fd_sc_hd__mux2_1 _4655_ (.A0(\core_0.execute.alu_mul_div.div_cur[13] ),
    .A1(_1513_),
    .S(_1409_),
    .X(_1514_));
 sky130_fd_sc_hd__or2_1 _4656_ (.A(_1415_),
    .B(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__o211a_1 _4657_ (.A1(\core_0.execute.alu_mul_div.div_cur[14] ),
    .A2(_1413_),
    .B1(_1515_),
    .C1(_1474_),
    .X(_0184_));
 sky130_fd_sc_hd__nand2_2 _4658_ (.A(_1409_),
    .B(_1412_),
    .Y(_1516_));
 sky130_fd_sc_hd__clkinv_2 _4659_ (.A(_1327_),
    .Y(_1517_));
 sky130_fd_sc_hd__or2_1 _4660_ (.A(_1517_),
    .B(_1408_),
    .X(_1518_));
 sky130_fd_sc_hd__xnor2_1 _4661_ (.A(_1407_),
    .B(_1518_),
    .Y(_1519_));
 sky130_fd_sc_hd__or2_1 _4662_ (.A(_1439_),
    .B(_1512_),
    .X(_1520_));
 sky130_fd_sc_hd__o211a_1 _4663_ (.A1(_1210_),
    .A2(_1519_),
    .B1(_1520_),
    .C1(_1410_),
    .X(_1521_));
 sky130_fd_sc_hd__a211o_1 _4664_ (.A1(\core_0.execute.alu_mul_div.div_cur[14] ),
    .A2(_1516_),
    .B1(_1416_),
    .C1(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__o211a_1 _4665_ (.A1(\core_0.execute.alu_mul_div.div_cur[15] ),
    .A2(_1413_),
    .B1(_1522_),
    .C1(_1474_),
    .X(_0185_));
 sky130_fd_sc_hd__or3_1 _4666_ (.A(\core_0.dec_l_reg_sel[2] ),
    .B(\core_0.dec_l_reg_sel[1] ),
    .C(_0709_),
    .X(_1523_));
 sky130_fd_sc_hd__buf_6 _4667_ (.A(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__nor2_4 _4668_ (.A(_0699_),
    .B(_0708_),
    .Y(_1525_));
 sky130_fd_sc_hd__buf_4 _4669_ (.A(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__and3b_4 _4670_ (.A_N(_0701_),
    .B(_0702_),
    .C(_0699_),
    .X(_1527_));
 sky130_fd_sc_hd__buf_2 _4671_ (.A(\core_0.dec_l_reg_sel[2] ),
    .X(_1528_));
 sky130_fd_sc_hd__buf_2 _4672_ (.A(\core_0.dec_l_reg_sel[1] ),
    .X(_1529_));
 sky130_fd_sc_hd__nor3b_2 _4673_ (.A(_1528_),
    .B(_0709_),
    .C_N(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__buf_4 _4674_ (.A(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__a22o_1 _4675_ (.A1(\core_0.execute.rf.reg_outputs[5][15] ),
    .A2(_1527_),
    .B1(_1531_),
    .B2(\core_0.execute.rf.reg_outputs[2][15] ),
    .X(_1532_));
 sky130_fd_sc_hd__a31o_1 _4676_ (.A1(\core_0.execute.rf.reg_outputs[1][15] ),
    .A2(_0714_),
    .A3(_1526_),
    .B1(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__and3b_1 _4677_ (.A_N(_0709_),
    .B(_0708_),
    .C(_1528_),
    .X(_1534_));
 sky130_fd_sc_hd__buf_4 _4678_ (.A(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__and2b_1 _4679_ (.A_N(\core_0.dec_l_reg_sel[2] ),
    .B(_1529_),
    .X(_1536_));
 sky130_fd_sc_hd__clkbuf_4 _4680_ (.A(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__a32o_1 _4681_ (.A1(\core_0.execute.rf.reg_outputs[3][15] ),
    .A2(_0713_),
    .A3(_1537_),
    .B1(_0703_),
    .B2(\core_0.execute.rf.reg_outputs[7][15] ),
    .X(_1538_));
 sky130_fd_sc_hd__o21a_1 _4682_ (.A1(\core_0.execute.rf.reg_outputs[4][15] ),
    .A2(_0717_),
    .B1(_0711_),
    .X(_1539_));
 sky130_fd_sc_hd__a211o_1 _4683_ (.A1(\core_0.execute.rf.reg_outputs[6][15] ),
    .A2(_1535_),
    .B1(_1538_),
    .C1(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__o22ai_4 _4684_ (.A1(net94),
    .A2(_1524_),
    .B1(_1533_),
    .B2(_1540_),
    .Y(_1541_));
 sky130_fd_sc_hd__inv_4 _4685_ (.A(_1541_),
    .Y(_1542_));
 sky130_fd_sc_hd__nor2_1 _4686_ (.A(_1210_),
    .B(_1425_),
    .Y(_1543_));
 sky130_fd_sc_hd__a22o_1 _4687_ (.A1(\core_0.execute.rf.reg_outputs[5][9] ),
    .A2(_1527_),
    .B1(_1531_),
    .B2(\core_0.execute.rf.reg_outputs[2][9] ),
    .X(_1544_));
 sky130_fd_sc_hd__a31o_1 _4688_ (.A1(\core_0.execute.rf.reg_outputs[1][9] ),
    .A2(_0714_),
    .A3(_1526_),
    .B1(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__o21a_1 _4689_ (.A1(\core_0.execute.rf.reg_outputs[4][9] ),
    .A2(_0717_),
    .B1(_0711_),
    .X(_1546_));
 sky130_fd_sc_hd__a32o_1 _4690_ (.A1(\core_0.execute.rf.reg_outputs[3][9] ),
    .A2(_0713_),
    .A3(_1537_),
    .B1(_0703_),
    .B2(\core_0.execute.rf.reg_outputs[7][9] ),
    .X(_1547_));
 sky130_fd_sc_hd__a211o_1 _4691_ (.A1(\core_0.execute.rf.reg_outputs[6][9] ),
    .A2(_1535_),
    .B1(_1546_),
    .C1(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__o22a_4 _4692_ (.A1(net103),
    .A2(_1524_),
    .B1(_1545_),
    .B2(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__buf_6 _4693_ (.A(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__o21a_1 _4694_ (.A1(\core_0.execute.rf.reg_outputs[4][10] ),
    .A2(_0717_),
    .B1(_0711_),
    .X(_1551_));
 sky130_fd_sc_hd__a31o_1 _4695_ (.A1(\core_0.execute.rf.reg_outputs[1][10] ),
    .A2(_0714_),
    .A3(_1526_),
    .B1(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__and2_1 _4696_ (.A(\core_0.execute.rf.reg_outputs[2][10] ),
    .B(_1531_),
    .X(_1553_));
 sky130_fd_sc_hd__a22o_1 _4697_ (.A1(\core_0.execute.rf.reg_outputs[7][10] ),
    .A2(_0703_),
    .B1(_1535_),
    .B2(\core_0.execute.rf.reg_outputs[6][10] ),
    .X(_1554_));
 sky130_fd_sc_hd__and3_1 _4698_ (.A(\core_0.execute.rf.reg_outputs[3][10] ),
    .B(_0713_),
    .C(_1537_),
    .X(_1555_));
 sky130_fd_sc_hd__a211o_1 _4699_ (.A1(\core_0.execute.rf.reg_outputs[5][10] ),
    .A2(_1527_),
    .B1(_1554_),
    .C1(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__o32a_4 _4700_ (.A1(_1552_),
    .A2(_1553_),
    .A3(_1556_),
    .B1(_1524_),
    .B2(net89),
    .X(_1557_));
 sky130_fd_sc_hd__buf_6 _4701_ (.A(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__clkinv_4 _4702_ (.A(\core_0.execute.alu_mul_div.cbit[0] ),
    .Y(_1559_));
 sky130_fd_sc_hd__clkbuf_8 _4703_ (.A(_1559_),
    .X(_1560_));
 sky130_fd_sc_hd__mux2_1 _4704_ (.A0(_1550_),
    .A1(_1558_),
    .S(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__nor3_2 _4705_ (.A(_1528_),
    .B(_0708_),
    .C(_0709_),
    .Y(_1562_));
 sky130_fd_sc_hd__buf_6 _4706_ (.A(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__a22o_1 _4707_ (.A1(\core_0.execute.rf.reg_outputs[1][7] ),
    .A2(_1525_),
    .B1(_1535_),
    .B2(\core_0.execute.rf.reg_outputs[6][7] ),
    .X(_1564_));
 sky130_fd_sc_hd__a32o_1 _4708_ (.A1(\core_0.execute.rf.reg_outputs[4][7] ),
    .A2(_0706_),
    .A3(_0711_),
    .B1(_1531_),
    .B2(\core_0.execute.rf.reg_outputs[2][7] ),
    .X(_1565_));
 sky130_fd_sc_hd__o21a_2 _4709_ (.A1(_1564_),
    .A2(_1565_),
    .B1(_1524_),
    .X(_1566_));
 sky130_fd_sc_hd__and2b_2 _4710_ (.A_N(_1529_),
    .B(\core_0.dec_l_reg_sel[2] ),
    .X(_1567_));
 sky130_fd_sc_hd__and3_1 _4711_ (.A(\core_0.execute.rf.reg_outputs[7][7] ),
    .B(_0699_),
    .C(_0701_),
    .X(_1568_));
 sky130_fd_sc_hd__a221o_2 _4712_ (.A1(\core_0.execute.rf.reg_outputs[3][7] ),
    .A2(_1537_),
    .B1(_1567_),
    .B2(\core_0.execute.rf.reg_outputs[5][7] ),
    .C1(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__and2_1 _4713_ (.A(_0714_),
    .B(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__a211o_4 _4714_ (.A1(net101),
    .A2(_1563_),
    .B1(_1566_),
    .C1(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__buf_6 _4715_ (.A(_1524_),
    .X(_1572_));
 sky130_fd_sc_hd__and2_2 _4716_ (.A(\core_0.execute.rf.reg_outputs[2][8] ),
    .B(_1531_),
    .X(_1573_));
 sky130_fd_sc_hd__and3_1 _4717_ (.A(\core_0.execute.rf.reg_outputs[1][8] ),
    .B(_0713_),
    .C(_1525_),
    .X(_1574_));
 sky130_fd_sc_hd__o21a_1 _4718_ (.A1(\core_0.execute.rf.reg_outputs[4][8] ),
    .A2(_0717_),
    .B1(_0711_),
    .X(_1575_));
 sky130_fd_sc_hd__and4b_1 _4719_ (.A_N(_0706_),
    .B(_0701_),
    .C(_0702_),
    .D(\core_0.execute.rf.reg_outputs[3][8] ),
    .X(_1576_));
 sky130_fd_sc_hd__a221o_1 _4720_ (.A1(\core_0.execute.rf.reg_outputs[7][8] ),
    .A2(_0703_),
    .B1(_1535_),
    .B2(\core_0.execute.rf.reg_outputs[6][8] ),
    .C1(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__a2111o_2 _4721_ (.A1(\core_0.execute.rf.reg_outputs[5][8] ),
    .A2(_1527_),
    .B1(_1574_),
    .C1(_1575_),
    .D1(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__o22a_4 _4722_ (.A1(net102),
    .A2(_1572_),
    .B1(_1573_),
    .B2(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__mux2_1 _4723_ (.A0(_1571_),
    .A1(_1579_),
    .S(_1560_),
    .X(_1580_));
 sky130_fd_sc_hd__mux2_1 _4724_ (.A0(_1561_),
    .A1(_1580_),
    .S(_1206_),
    .X(_1581_));
 sky130_fd_sc_hd__and4bb_1 _4725_ (.A_N(_0706_),
    .B_N(_0704_),
    .C(_0713_),
    .D(\core_0.execute.rf.reg_outputs[1][12] ),
    .X(_1582_));
 sky130_fd_sc_hd__a221o_1 _4726_ (.A1(\core_0.execute.rf.reg_outputs[5][12] ),
    .A2(_1527_),
    .B1(_1531_),
    .B2(\core_0.execute.rf.reg_outputs[2][12] ),
    .C1(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__a32o_1 _4727_ (.A1(\core_0.execute.rf.reg_outputs[3][12] ),
    .A2(_0714_),
    .A3(_1537_),
    .B1(_0703_),
    .B2(\core_0.execute.rf.reg_outputs[7][12] ),
    .X(_1584_));
 sky130_fd_sc_hd__or2b_1 _4728_ (.A(\core_0.execute.rf.reg_outputs[4][12] ),
    .B_N(_0706_),
    .X(_1585_));
 sky130_fd_sc_hd__a22o_1 _4729_ (.A1(\core_0.execute.rf.reg_outputs[6][12] ),
    .A2(_1535_),
    .B1(_1585_),
    .B2(_0711_),
    .X(_1586_));
 sky130_fd_sc_hd__or3_2 _4730_ (.A(_1583_),
    .B(_1584_),
    .C(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__o21a_4 _4731_ (.A1(net91),
    .A2(_1572_),
    .B1(_1587_),
    .X(_1588_));
 sky130_fd_sc_hd__a22o_1 _4732_ (.A1(\core_0.execute.rf.reg_outputs[5][11] ),
    .A2(_1527_),
    .B1(_1531_),
    .B2(\core_0.execute.rf.reg_outputs[2][11] ),
    .X(_1589_));
 sky130_fd_sc_hd__a31o_2 _4733_ (.A1(\core_0.execute.rf.reg_outputs[1][11] ),
    .A2(_0714_),
    .A3(_1526_),
    .B1(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__or2_1 _4734_ (.A(\core_0.execute.rf.reg_outputs[4][11] ),
    .B(_0717_),
    .X(_1591_));
 sky130_fd_sc_hd__a32o_1 _4735_ (.A1(\core_0.execute.rf.reg_outputs[3][11] ),
    .A2(_0713_),
    .A3(_1537_),
    .B1(_0703_),
    .B2(\core_0.execute.rf.reg_outputs[7][11] ),
    .X(_1592_));
 sky130_fd_sc_hd__a221o_4 _4736_ (.A1(\core_0.execute.rf.reg_outputs[6][11] ),
    .A2(_1535_),
    .B1(_1591_),
    .B2(_0711_),
    .C1(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__o22a_4 _4737_ (.A1(net90),
    .A2(_1524_),
    .B1(_1590_),
    .B2(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__mux2_1 _4738_ (.A0(_1588_),
    .A1(_1594_),
    .S(_1205_),
    .X(_1595_));
 sky130_fd_sc_hd__a22o_1 _4739_ (.A1(\core_0.execute.rf.reg_outputs[2][13] ),
    .A2(_1531_),
    .B1(_1535_),
    .B2(\core_0.execute.rf.reg_outputs[6][13] ),
    .X(_1596_));
 sky130_fd_sc_hd__a31o_2 _4740_ (.A1(\core_0.execute.rf.reg_outputs[3][13] ),
    .A2(_0715_),
    .A3(_1537_),
    .B1(_1596_),
    .X(_1597_));
 sky130_fd_sc_hd__or2b_1 _4741_ (.A(\core_0.execute.rf.reg_outputs[4][13] ),
    .B_N(_0706_),
    .X(_1598_));
 sky130_fd_sc_hd__a32o_1 _4742_ (.A1(\core_0.execute.rf.reg_outputs[1][13] ),
    .A2(_0714_),
    .A3(_1526_),
    .B1(_1598_),
    .B2(_0711_),
    .X(_1599_));
 sky130_fd_sc_hd__a221o_2 _4743_ (.A1(\core_0.execute.rf.reg_outputs[7][13] ),
    .A2(_0703_),
    .B1(_1527_),
    .B2(\core_0.execute.rf.reg_outputs[5][13] ),
    .C1(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__o22a_4 _4744_ (.A1(net92),
    .A2(_1572_),
    .B1(_1597_),
    .B2(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__nor2_8 _4745_ (.A(_1560_),
    .B(_1207_),
    .Y(_1602_));
 sky130_fd_sc_hd__or2_1 _4746_ (.A(_1205_),
    .B(_1207_),
    .X(_1603_));
 sky130_fd_sc_hd__a22o_2 _4747_ (.A1(\core_0.execute.rf.reg_outputs[7][14] ),
    .A2(_0703_),
    .B1(_1535_),
    .B2(\core_0.execute.rf.reg_outputs[6][14] ),
    .X(_1604_));
 sky130_fd_sc_hd__and3_1 _4748_ (.A(\core_0.execute.rf.reg_outputs[3][14] ),
    .B(_0713_),
    .C(_1537_),
    .X(_1605_));
 sky130_fd_sc_hd__o21a_1 _4749_ (.A1(\core_0.execute.rf.reg_outputs[4][14] ),
    .A2(_0717_),
    .B1(_0711_),
    .X(_1606_));
 sky130_fd_sc_hd__a32o_1 _4750_ (.A1(\core_0.execute.rf.reg_outputs[1][14] ),
    .A2(_0714_),
    .A3(_1526_),
    .B1(_1527_),
    .B2(\core_0.execute.rf.reg_outputs[5][14] ),
    .X(_1607_));
 sky130_fd_sc_hd__a2111o_2 _4751_ (.A1(\core_0.execute.rf.reg_outputs[2][14] ),
    .A2(_1531_),
    .B1(_1605_),
    .C1(_1606_),
    .D1(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__o22ai_4 _4752_ (.A1(net93),
    .A2(_1572_),
    .B1(_1604_),
    .B2(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__nor2_1 _4753_ (.A(_1603_),
    .B(_1609_),
    .Y(_1610_));
 sky130_fd_sc_hd__a221o_1 _4754_ (.A1(_1207_),
    .A2(_1595_),
    .B1(_1601_),
    .B2(_1602_),
    .C1(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__mux2_1 _4755_ (.A0(_1581_),
    .A1(_1611_),
    .S(_1204_),
    .X(_1612_));
 sky130_fd_sc_hd__or4bb_1 _4756_ (.A(_1529_),
    .B(_0709_),
    .C_N(\core_0.execute.rf.reg_outputs[4][1] ),
    .D_N(_1528_),
    .X(_1613_));
 sky130_fd_sc_hd__or3b_1 _4757_ (.A(_1528_),
    .B(_1529_),
    .C_N(\core_0.execute.rf.reg_outputs[1][1] ),
    .X(_1614_));
 sky130_fd_sc_hd__nand4b_1 _4758_ (.A_N(_0702_),
    .B(_0708_),
    .C(_0699_),
    .D(\core_0.execute.rf.reg_outputs[6][1] ),
    .Y(_1615_));
 sky130_fd_sc_hd__or4bb_1 _4759_ (.A(_1528_),
    .B(_0709_),
    .C_N(_1529_),
    .D_N(\core_0.execute.rf.reg_outputs[2][1] ),
    .X(_1616_));
 sky130_fd_sc_hd__a41o_1 _4760_ (.A1(_1613_),
    .A2(_1614_),
    .A3(_1615_),
    .A4(_1616_),
    .B1(_1562_),
    .X(_1617_));
 sky130_fd_sc_hd__nand3_2 _4761_ (.A(\core_0.execute.rf.reg_outputs[7][1] ),
    .B(_0699_),
    .C(_0708_),
    .Y(_1618_));
 sky130_fd_sc_hd__nand3b_2 _4762_ (.A_N(_0708_),
    .B(_0699_),
    .C(\core_0.execute.rf.reg_outputs[5][1] ),
    .Y(_1619_));
 sky130_fd_sc_hd__nand3b_2 _4763_ (.A_N(_0699_),
    .B(_0708_),
    .C(\core_0.execute.rf.reg_outputs[3][1] ),
    .Y(_1620_));
 sky130_fd_sc_hd__a31o_1 _4764_ (.A1(_1618_),
    .A2(_1619_),
    .A3(_1620_),
    .B1(_0705_),
    .X(_1621_));
 sky130_fd_sc_hd__nand2_1 _4765_ (.A(net95),
    .B(_1562_),
    .Y(_1622_));
 sky130_fd_sc_hd__and3_1 _4766_ (.A(_1617_),
    .B(_1621_),
    .C(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__buf_4 _4767_ (.A(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__and3_1 _4768_ (.A(\core_0.execute.rf.reg_outputs[7][2] ),
    .B(_0700_),
    .C(_0701_),
    .X(_1625_));
 sky130_fd_sc_hd__a221o_4 _4769_ (.A1(\core_0.execute.rf.reg_outputs[3][2] ),
    .A2(_1537_),
    .B1(_1567_),
    .B2(\core_0.execute.rf.reg_outputs[5][2] ),
    .C1(_1625_),
    .X(_1626_));
 sky130_fd_sc_hd__and4bb_1 _4770_ (.A_N(_0700_),
    .B_N(_0702_),
    .C(_0701_),
    .D(\core_0.execute.rf.reg_outputs[2][2] ),
    .X(_1627_));
 sky130_fd_sc_hd__and4bb_1 _4771_ (.A_N(_0701_),
    .B_N(_0702_),
    .C(\core_0.execute.rf.reg_outputs[4][2] ),
    .D(_0700_),
    .X(_1628_));
 sky130_fd_sc_hd__and4b_1 _4772_ (.A_N(_0702_),
    .B(_0701_),
    .C(_0700_),
    .D(\core_0.execute.rf.reg_outputs[6][2] ),
    .X(_1629_));
 sky130_fd_sc_hd__nor3b_4 _4773_ (.A(_0706_),
    .B(_0704_),
    .C_N(\core_0.execute.rf.reg_outputs[1][2] ),
    .Y(_1630_));
 sky130_fd_sc_hd__o41a_2 _4774_ (.A1(_1627_),
    .A2(_1628_),
    .A3(_1629_),
    .A4(_1630_),
    .B1(_1524_),
    .X(_1631_));
 sky130_fd_sc_hd__a221oi_4 _4775_ (.A1(net96),
    .A2(_1563_),
    .B1(_1626_),
    .B2(_0715_),
    .C1(_1631_),
    .Y(_1632_));
 sky130_fd_sc_hd__clkbuf_4 _4776_ (.A(_1632_),
    .X(_1633_));
 sky130_fd_sc_hd__mux2_1 _4777_ (.A0(_1624_),
    .A1(_1633_),
    .S(_1559_),
    .X(_1634_));
 sky130_fd_sc_hd__and4b_1 _4778_ (.A_N(_0709_),
    .B(\core_0.dec_l_reg_sel[1] ),
    .C(\core_0.dec_l_reg_sel[2] ),
    .D(\core_0.execute.rf.reg_outputs[6][0] ),
    .X(_1635_));
 sky130_fd_sc_hd__nor3b_1 _4779_ (.A(_1528_),
    .B(_1529_),
    .C_N(\core_0.execute.rf.reg_outputs[1][0] ),
    .Y(_1636_));
 sky130_fd_sc_hd__and4bb_1 _4780_ (.A_N(\core_0.dec_l_reg_sel[2] ),
    .B_N(_0709_),
    .C(\core_0.dec_l_reg_sel[1] ),
    .D(\core_0.execute.rf.reg_outputs[2][0] ),
    .X(_1637_));
 sky130_fd_sc_hd__and4bb_1 _4781_ (.A_N(\core_0.dec_l_reg_sel[1] ),
    .B_N(_0709_),
    .C(\core_0.execute.rf.reg_outputs[4][0] ),
    .D(\core_0.dec_l_reg_sel[2] ),
    .X(_1638_));
 sky130_fd_sc_hd__o41a_2 _4782_ (.A1(_1635_),
    .A2(_1636_),
    .A3(_1637_),
    .A4(_1638_),
    .B1(_1523_),
    .X(_1639_));
 sky130_fd_sc_hd__and3_1 _4783_ (.A(\core_0.execute.rf.reg_outputs[7][0] ),
    .B(\core_0.dec_l_reg_sel[2] ),
    .C(\core_0.dec_l_reg_sel[1] ),
    .X(_1640_));
 sky130_fd_sc_hd__and3b_1 _4784_ (.A_N(_1529_),
    .B(\core_0.dec_l_reg_sel[2] ),
    .C(\core_0.execute.rf.reg_outputs[5][0] ),
    .X(_1641_));
 sky130_fd_sc_hd__and3b_1 _4785_ (.A_N(_1528_),
    .B(_1529_),
    .C(\core_0.execute.rf.reg_outputs[3][0] ),
    .X(_1642_));
 sky130_fd_sc_hd__o31a_1 _4786_ (.A1(_1640_),
    .A2(_1641_),
    .A3(_1642_),
    .B1(_0702_),
    .X(_1643_));
 sky130_fd_sc_hd__a211o_4 _4787_ (.A1(net88),
    .A2(_1562_),
    .B1(_1639_),
    .C1(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__and2_2 _4788_ (.A(_1559_),
    .B(\core_0.execute.alu_mul_div.cbit[1] ),
    .X(_1645_));
 sky130_fd_sc_hd__a2bb2o_2 _4789_ (.A1_N(_1206_),
    .A2_N(_1634_),
    .B1(_1644_),
    .B2(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__clkinv_2 _4790_ (.A(_1646_),
    .Y(_1647_));
 sky130_fd_sc_hd__and3_1 _4791_ (.A(\core_0.execute.rf.reg_outputs[7][6] ),
    .B(_1528_),
    .C(_0708_),
    .X(_1648_));
 sky130_fd_sc_hd__a221o_2 _4792_ (.A1(\core_0.execute.rf.reg_outputs[3][6] ),
    .A2(_1536_),
    .B1(_1567_),
    .B2(\core_0.execute.rf.reg_outputs[5][6] ),
    .C1(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__and2_1 _4793_ (.A(_0713_),
    .B(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__a32o_1 _4794_ (.A1(\core_0.execute.rf.reg_outputs[4][6] ),
    .A2(_0700_),
    .A3(_0710_),
    .B1(_1525_),
    .B2(\core_0.execute.rf.reg_outputs[1][6] ),
    .X(_1651_));
 sky130_fd_sc_hd__or2_1 _4795_ (.A(_1563_),
    .B(_1651_),
    .X(_1652_));
 sky130_fd_sc_hd__a22o_2 _4796_ (.A1(\core_0.execute.rf.reg_outputs[2][6] ),
    .A2(_1531_),
    .B1(_1535_),
    .B2(\core_0.execute.rf.reg_outputs[6][6] ),
    .X(_1653_));
 sky130_fd_sc_hd__o32a_4 _4797_ (.A1(_1650_),
    .A2(_1652_),
    .A3(_1653_),
    .B1(_1524_),
    .B2(net100),
    .X(_1654_));
 sky130_fd_sc_hd__a22o_1 _4798_ (.A1(\core_0.execute.rf.reg_outputs[1][5] ),
    .A2(_1525_),
    .B1(_1534_),
    .B2(\core_0.execute.rf.reg_outputs[6][5] ),
    .X(_1655_));
 sky130_fd_sc_hd__a32o_1 _4799_ (.A1(\core_0.execute.rf.reg_outputs[4][5] ),
    .A2(_0700_),
    .A3(_0710_),
    .B1(_1530_),
    .B2(\core_0.execute.rf.reg_outputs[2][5] ),
    .X(_1656_));
 sky130_fd_sc_hd__o21a_2 _4800_ (.A1(_1655_),
    .A2(_1656_),
    .B1(_1523_),
    .X(_1657_));
 sky130_fd_sc_hd__and3_1 _4801_ (.A(\core_0.execute.rf.reg_outputs[7][5] ),
    .B(_0699_),
    .C(_0708_),
    .X(_1658_));
 sky130_fd_sc_hd__a221o_2 _4802_ (.A1(\core_0.execute.rf.reg_outputs[3][5] ),
    .A2(_1536_),
    .B1(_1567_),
    .B2(\core_0.execute.rf.reg_outputs[5][5] ),
    .C1(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__and2_1 _4803_ (.A(_0714_),
    .B(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__a211o_4 _4804_ (.A1(net99),
    .A2(_1563_),
    .B1(_1657_),
    .C1(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__mux2_1 _4805_ (.A0(_1654_),
    .A1(_1661_),
    .S(_1205_),
    .X(_1662_));
 sky130_fd_sc_hd__clkinv_2 _4806_ (.A(_1662_),
    .Y(_1663_));
 sky130_fd_sc_hd__and3_1 _4807_ (.A(\core_0.execute.rf.reg_outputs[7][3] ),
    .B(_0700_),
    .C(_0701_),
    .X(_1664_));
 sky130_fd_sc_hd__a221o_4 _4808_ (.A1(\core_0.execute.rf.reg_outputs[3][3] ),
    .A2(_1537_),
    .B1(_1567_),
    .B2(\core_0.execute.rf.reg_outputs[5][3] ),
    .C1(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__and2_1 _4809_ (.A(\core_0.execute.rf.reg_outputs[6][3] ),
    .B(_1534_),
    .X(_1666_));
 sky130_fd_sc_hd__and2_1 _4810_ (.A(\core_0.execute.rf.reg_outputs[1][3] ),
    .B(_1525_),
    .X(_1667_));
 sky130_fd_sc_hd__a32o_1 _4811_ (.A1(\core_0.execute.rf.reg_outputs[4][3] ),
    .A2(_0706_),
    .A3(_0710_),
    .B1(_1530_),
    .B2(\core_0.execute.rf.reg_outputs[2][3] ),
    .X(_1668_));
 sky130_fd_sc_hd__o31a_1 _4812_ (.A1(_1666_),
    .A2(_1667_),
    .A3(_1668_),
    .B1(_1524_),
    .X(_1669_));
 sky130_fd_sc_hd__a221oi_4 _4813_ (.A1(net97),
    .A2(_1563_),
    .B1(_1665_),
    .B2(_0715_),
    .C1(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__a32o_1 _4814_ (.A1(\core_0.execute.rf.reg_outputs[4][4] ),
    .A2(_0699_),
    .A3(_0710_),
    .B1(_1530_),
    .B2(\core_0.execute.rf.reg_outputs[2][4] ),
    .X(_1671_));
 sky130_fd_sc_hd__a221o_1 _4815_ (.A1(\core_0.execute.rf.reg_outputs[1][4] ),
    .A2(_1525_),
    .B1(_1534_),
    .B2(\core_0.execute.rf.reg_outputs[6][4] ),
    .C1(_1671_),
    .X(_1672_));
 sky130_fd_sc_hd__and3_1 _4816_ (.A(\core_0.execute.rf.reg_outputs[7][4] ),
    .B(_1528_),
    .C(_1529_),
    .X(_1673_));
 sky130_fd_sc_hd__a221o_2 _4817_ (.A1(\core_0.execute.rf.reg_outputs[3][4] ),
    .A2(_1536_),
    .B1(_1567_),
    .B2(\core_0.execute.rf.reg_outputs[5][4] ),
    .C1(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__a22o_1 _4818_ (.A1(net98),
    .A2(_1563_),
    .B1(_1674_),
    .B2(_0713_),
    .X(_1675_));
 sky130_fd_sc_hd__a21oi_2 _4819_ (.A1(_1524_),
    .A2(_1672_),
    .B1(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__buf_4 _4820_ (.A(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__mux2_1 _4821_ (.A0(_1670_),
    .A1(_1677_),
    .S(_1560_),
    .X(_1678_));
 sky130_fd_sc_hd__mux2_1 _4822_ (.A0(_1663_),
    .A1(_1678_),
    .S(_1206_),
    .X(_1679_));
 sky130_fd_sc_hd__mux2_1 _4823_ (.A0(_1647_),
    .A1(_1679_),
    .S(_1204_),
    .X(_1680_));
 sky130_fd_sc_hd__inv_2 _4824_ (.A(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__mux2_1 _4825_ (.A0(_1612_),
    .A1(_1681_),
    .S(_1202_),
    .X(_1682_));
 sky130_fd_sc_hd__or3_1 _4826_ (.A(_1415_),
    .B(_1543_),
    .C(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__o211a_1 _4827_ (.A1(\core_0.execute.alu_mul_div.div_cur[0] ),
    .A2(_1413_),
    .B1(_1683_),
    .C1(_0742_),
    .X(_1684_));
 sky130_fd_sc_hd__a31o_1 _4828_ (.A1(\core_0.decode.o_submit ),
    .A2(_1411_),
    .A3(_1542_),
    .B1(_1684_),
    .X(_0186_));
 sky130_fd_sc_hd__a21oi_1 _4829_ (.A1(\core_0.dec_jump_cond_code[4] ),
    .A2(_1062_),
    .B1(\core_0.dec_pc_inc ),
    .Y(_1685_));
 sky130_fd_sc_hd__and2b_1 _4830_ (.A_N(_1685_),
    .B(_0746_),
    .X(_1686_));
 sky130_fd_sc_hd__buf_4 _4831_ (.A(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__or2_1 _4832_ (.A(net72),
    .B(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__inv_2 _4833_ (.A(_1062_),
    .Y(_1689_));
 sky130_fd_sc_hd__a21o_1 _4834_ (.A1(\core_0.dec_jump_cond_code[4] ),
    .A2(_1689_),
    .B1(_1039_),
    .X(_1690_));
 sky130_fd_sc_hd__nand2_4 _4835_ (.A(_0746_),
    .B(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__clkbuf_4 _4836_ (.A(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__nand2_1 _4837_ (.A(net72),
    .B(_1687_),
    .Y(_1693_));
 sky130_fd_sc_hd__a31o_1 _4838_ (.A1(_1688_),
    .A2(_1692_),
    .A3(_1693_),
    .B1(_0674_),
    .X(_1694_));
 sky130_fd_sc_hd__or2_1 _4839_ (.A(_1038_),
    .B(_1152_),
    .X(_1695_));
 sky130_fd_sc_hd__clkinv_2 _4840_ (.A(\core_0.execute.alu_mul_div.i_mod ),
    .Y(_1696_));
 sky130_fd_sc_hd__clkbuf_4 _4841_ (.A(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__o21a_4 _4842_ (.A1(_1077_),
    .A2(_0647_),
    .B1(_1373_),
    .X(_1698_));
 sky130_fd_sc_hd__nand4_2 _4843_ (.A(_1379_),
    .B(_1380_),
    .C(_1376_),
    .D(_1377_),
    .Y(_1699_));
 sky130_fd_sc_hd__nor2_2 _4844_ (.A(_1698_),
    .B(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__o21ai_4 _4845_ (.A1(_1077_),
    .A2(_0633_),
    .B1(_1364_),
    .Y(_1701_));
 sky130_fd_sc_hd__inv_2 _4846_ (.A(\core_0.decode.oc_alu_mode[12] ),
    .Y(_1702_));
 sky130_fd_sc_hd__mux2_4 _4847_ (.A0(net187),
    .A1(net203),
    .S(_1341_),
    .X(_1703_));
 sky130_fd_sc_hd__or4_1 _4848_ (.A(_1702_),
    .B(_1703_),
    .C(_1698_),
    .D(_1699_),
    .X(_1704_));
 sky130_fd_sc_hd__xnor2_2 _4849_ (.A(_1701_),
    .B(_1704_),
    .Y(_1705_));
 sky130_fd_sc_hd__o21ai_1 _4850_ (.A1(\core_0.decode.oc_alu_mode[12] ),
    .A2(\core_0.decode.oc_alu_mode[13] ),
    .B1(_1362_),
    .Y(_1706_));
 sky130_fd_sc_hd__nor2_4 _4851_ (.A(_1705_),
    .B(_1706_),
    .Y(_1707_));
 sky130_fd_sc_hd__nor2_1 _4852_ (.A(\core_0.decode.oc_alu_mode[12] ),
    .B(_1644_),
    .Y(_1708_));
 sky130_fd_sc_hd__a21oi_4 _4853_ (.A1(_1341_),
    .A2(_0627_),
    .B1(_1361_),
    .Y(_1709_));
 sky130_fd_sc_hd__a2111o_1 _4854_ (.A1(_1076_),
    .A2(net191),
    .B1(_1352_),
    .C1(_1355_),
    .D1(_1356_),
    .X(_1710_));
 sky130_fd_sc_hd__or4_1 _4855_ (.A(_1323_),
    .B(_1325_),
    .C(_1328_),
    .D(_1330_),
    .X(_1711_));
 sky130_fd_sc_hd__a2111o_1 _4856_ (.A1(_1077_),
    .A2(net182),
    .B1(_1333_),
    .C1(_1336_),
    .D1(_1337_),
    .X(_1712_));
 sky130_fd_sc_hd__o41a_1 _4857_ (.A1(_1709_),
    .A2(_1710_),
    .A3(_1711_),
    .A4(_1712_),
    .B1(\core_0.decode.oc_alu_mode[12] ),
    .X(_1713_));
 sky130_fd_sc_hd__o311a_1 _4858_ (.A1(_1703_),
    .A2(_1698_),
    .A3(_1699_),
    .B1(_1701_),
    .C1(\core_0.decode.oc_alu_mode[12] ),
    .X(_1714_));
 sky130_fd_sc_hd__or4_2 _4859_ (.A(_1493_),
    .B(_1344_),
    .C(_1482_),
    .D(_1391_),
    .X(_1715_));
 sky130_fd_sc_hd__a211o_1 _4860_ (.A1(_1341_),
    .A2(_0627_),
    .B1(_1361_),
    .C1(_1702_),
    .X(_1716_));
 sky130_fd_sc_hd__a211o_1 _4861_ (.A1(_1710_),
    .A2(_1716_),
    .B1(_1712_),
    .C1(_1711_),
    .X(_1717_));
 sky130_fd_sc_hd__or4_2 _4862_ (.A(_1713_),
    .B(_1714_),
    .C(_1715_),
    .D(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__buf_2 _4863_ (.A(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__nor2_1 _4864_ (.A(_1702_),
    .B(_1542_),
    .Y(_1720_));
 sky130_fd_sc_hd__buf_2 _4865_ (.A(_1720_),
    .X(_1721_));
 sky130_fd_sc_hd__nor2_2 _4866_ (.A(_1719_),
    .B(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__and2b_1 _4867_ (.A_N(_1708_),
    .B(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__nand2_2 _4868_ (.A(_1379_),
    .B(_1380_),
    .Y(_1724_));
 sky130_fd_sc_hd__buf_4 _4869_ (.A(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__or4_1 _4870_ (.A(_1709_),
    .B(_1710_),
    .C(_1711_),
    .D(_1712_),
    .X(_1726_));
 sky130_fd_sc_hd__or2_1 _4871_ (.A(_1726_),
    .B(_1715_),
    .X(_1727_));
 sky130_fd_sc_hd__clkbuf_4 _4872_ (.A(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__nand2_4 _4873_ (.A(_1376_),
    .B(_1377_),
    .Y(_1729_));
 sky130_fd_sc_hd__mux2_1 _4874_ (.A0(_1633_),
    .A1(_1670_),
    .S(_1729_),
    .X(_1730_));
 sky130_fd_sc_hd__nor2_1 _4875_ (.A(_1728_),
    .B(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__clkinv_2 _4876_ (.A(_1624_),
    .Y(_1732_));
 sky130_fd_sc_hd__buf_2 _4877_ (.A(_1726_),
    .X(_1733_));
 sky130_fd_sc_hd__clkbuf_4 _4878_ (.A(_1715_),
    .X(_1734_));
 sky130_fd_sc_hd__nor2_1 _4879_ (.A(_1733_),
    .B(_1734_),
    .Y(_1735_));
 sky130_fd_sc_hd__or3_2 _4880_ (.A(_1419_),
    .B(_1420_),
    .C(_1644_),
    .X(_1736_));
 sky130_fd_sc_hd__and2_1 _4881_ (.A(_1379_),
    .B(_1380_),
    .X(_1737_));
 sky130_fd_sc_hd__buf_4 _4882_ (.A(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__buf_4 _4883_ (.A(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__o2111a_1 _4884_ (.A1(_1422_),
    .A2(_1732_),
    .B1(_1735_),
    .C1(_1736_),
    .D1(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__clkbuf_4 _4885_ (.A(_1698_),
    .X(_1741_));
 sky130_fd_sc_hd__a211o_1 _4886_ (.A1(_1725_),
    .A2(_1731_),
    .B1(_1740_),
    .C1(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__a211oi_4 _4887_ (.A1(net99),
    .A2(_1563_),
    .B1(_1657_),
    .C1(_1660_),
    .Y(_1743_));
 sky130_fd_sc_hd__mux2_1 _4888_ (.A0(_1743_),
    .A1(_1677_),
    .S(_1421_),
    .X(_1744_));
 sky130_fd_sc_hd__a211oi_4 _4889_ (.A1(net101),
    .A2(_1563_),
    .B1(_1566_),
    .C1(_1570_),
    .Y(_1745_));
 sky130_fd_sc_hd__o32ai_4 _4890_ (.A1(_1650_),
    .A2(_1652_),
    .A3(_1653_),
    .B1(_1572_),
    .B2(net100),
    .Y(_1746_));
 sky130_fd_sc_hd__mux2_1 _4891_ (.A0(_1745_),
    .A1(_1746_),
    .S(_1421_),
    .X(_1747_));
 sky130_fd_sc_hd__mux2_1 _4892_ (.A0(_1744_),
    .A1(_1747_),
    .S(_1725_),
    .X(_1748_));
 sky130_fd_sc_hd__buf_6 _4893_ (.A(_1741_),
    .X(_1749_));
 sky130_fd_sc_hd__o21ai_1 _4894_ (.A1(_1728_),
    .A2(_1748_),
    .B1(_1749_),
    .Y(_1750_));
 sky130_fd_sc_hd__buf_4 _4895_ (.A(_1703_),
    .X(_1751_));
 sky130_fd_sc_hd__nor2_1 _4896_ (.A(\core_0.decode.oc_alu_mode[1] ),
    .B(\core_0.decode.oc_alu_mode[12] ),
    .Y(_1752_));
 sky130_fd_sc_hd__or2_2 _4897_ (.A(_1701_),
    .B(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__nor2_2 _4898_ (.A(_1751_),
    .B(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__mux2_1 _4899_ (.A0(_1541_),
    .A1(_1609_),
    .S(_1421_),
    .X(_1755_));
 sky130_fd_sc_hd__o21ai_4 _4900_ (.A1(net91),
    .A2(_1572_),
    .B1(_1587_),
    .Y(_1756_));
 sky130_fd_sc_hd__o22ai_4 _4901_ (.A1(net92),
    .A2(_1572_),
    .B1(_1597_),
    .B2(_1600_),
    .Y(_1757_));
 sky130_fd_sc_hd__mux2_1 _4902_ (.A0(_1756_),
    .A1(_1757_),
    .S(_1729_),
    .X(_1758_));
 sky130_fd_sc_hd__mux2_1 _4903_ (.A0(_1755_),
    .A1(_1758_),
    .S(_1738_),
    .X(_1759_));
 sky130_fd_sc_hd__mux4_1 _4904_ (.A0(_1550_),
    .A1(_1579_),
    .A2(_1594_),
    .A3(_1558_),
    .S0(_1421_),
    .S1(_1724_),
    .X(_1760_));
 sky130_fd_sc_hd__nor2_1 _4905_ (.A(_1698_),
    .B(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__a2111oi_4 _4906_ (.A1(_1741_),
    .A2(_1759_),
    .B1(_1761_),
    .C1(_1728_),
    .D1(_1753_),
    .Y(_1762_));
 sky130_fd_sc_hd__and2_2 _4907_ (.A(\core_0.execute.alu_flag_reg.o_d[1] ),
    .B(\core_0.dec_alu_carry_en ),
    .X(_1763_));
 sky130_fd_sc_hd__buf_4 _4908_ (.A(_1729_),
    .X(_1764_));
 sky130_fd_sc_hd__nor2_1 _4909_ (.A(_1764_),
    .B(_1644_),
    .Y(_1765_));
 sky130_fd_sc_hd__a211oi_4 _4910_ (.A1(net88),
    .A2(_1563_),
    .B1(_1639_),
    .C1(_1643_),
    .Y(_1766_));
 sky130_fd_sc_hd__a21oi_4 _4911_ (.A1(_1376_),
    .A2(_1377_),
    .B1(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__nor2_1 _4912_ (.A(_1765_),
    .B(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__nand2_1 _4913_ (.A(_1763_),
    .B(_1768_),
    .Y(_1769_));
 sky130_fd_sc_hd__o22a_1 _4914_ (.A1(\core_0.decode.oc_alu_mode[4] ),
    .A2(\core_0.decode.oc_alu_mode[11] ),
    .B1(_1763_),
    .B2(_1768_),
    .X(_1770_));
 sky130_fd_sc_hd__or4_1 _4915_ (.A(\core_0.decode.oc_alu_mode[9] ),
    .B(\core_0.decode.oc_alu_mode[13] ),
    .C(\core_0.decode.oc_alu_mode[3] ),
    .D(\core_0.decode.oc_alu_mode[2] ),
    .X(_1771_));
 sky130_fd_sc_hd__or4_1 _4916_ (.A(\core_0.decode.oc_alu_mode[1] ),
    .B(\core_0.decode.oc_alu_mode[6] ),
    .C(\core_0.decode.oc_alu_mode[7] ),
    .D(\core_0.decode.oc_alu_mode[12] ),
    .X(_1772_));
 sky130_fd_sc_hd__inv_2 _4917_ (.A(\core_0.decode.oc_alu_mode[4] ),
    .Y(_1773_));
 sky130_fd_sc_hd__inv_4 _4918_ (.A(\core_0.decode.oc_alu_mode[11] ),
    .Y(_1774_));
 sky130_fd_sc_hd__and4bb_4 _4919_ (.A_N(_1771_),
    .B_N(_1772_),
    .C(_1773_),
    .D(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__or2_2 _4920_ (.A(\core_0.decode.oc_alu_mode[3] ),
    .B(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__a22o_1 _4921_ (.A1(\core_0.decode.oc_alu_mode[7] ),
    .A2(_1729_),
    .B1(_1644_),
    .B2(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__a21o_1 _4922_ (.A1(\core_0.decode.oc_alu_mode[9] ),
    .A2(_1736_),
    .B1(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__a221o_1 _4923_ (.A1(\core_0.decode.oc_alu_mode[2] ),
    .A2(_1767_),
    .B1(_1768_),
    .B2(\core_0.decode.oc_alu_mode[6] ),
    .C1(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__a221o_1 _4924_ (.A1(_1751_),
    .A2(_1762_),
    .B1(_1769_),
    .B2(_1770_),
    .C1(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__a31o_1 _4925_ (.A1(_1742_),
    .A2(_1750_),
    .A3(_1754_),
    .B1(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__a41o_2 _4926_ (.A1(_1371_),
    .A2(_1700_),
    .A3(_1707_),
    .A4(_1723_),
    .B1(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__or2_1 _4927_ (.A(\core_0.execute.alu_mul_div.i_mul ),
    .B(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__inv_2 _4928_ (.A(\core_0.execute.alu_mul_div.i_mul ),
    .Y(_1784_));
 sky130_fd_sc_hd__o21ba_1 _4929_ (.A1(_1784_),
    .A2(\core_0.execute.alu_mul_div.mul_res[0] ),
    .B1_N(_0988_),
    .X(_1785_));
 sky130_fd_sc_hd__a221o_1 _4930_ (.A1(\core_0.execute.alu_mul_div.div_res[0] ),
    .A2(_0989_),
    .B1(_1783_),
    .B2(_1785_),
    .C1(\core_0.execute.alu_mul_div.i_mod ),
    .X(_1786_));
 sky130_fd_sc_hd__o21a_2 _4931_ (.A1(_1697_),
    .A2(\core_0.execute.alu_mul_div.div_cur[0] ),
    .B1(_1786_),
    .X(_1787_));
 sky130_fd_sc_hd__clkinv_4 _4932_ (.A(\core_0.dec_sreg_irt ),
    .Y(_1788_));
 sky130_fd_sc_hd__buf_4 _4933_ (.A(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__nand2_2 _4934_ (.A(_1789_),
    .B(_1152_),
    .Y(_1790_));
 sky130_fd_sc_hd__buf_2 _4935_ (.A(_1691_),
    .X(_1791_));
 sky130_fd_sc_hd__nor2_2 _4936_ (.A(\core_0.execute.sreg_irq_pc.o_d[0] ),
    .B(_1788_),
    .Y(_1792_));
 sky130_fd_sc_hd__nor2_1 _4937_ (.A(_1791_),
    .B(_1792_),
    .Y(_1793_));
 sky130_fd_sc_hd__o221a_1 _4938_ (.A1(_1695_),
    .A2(_1787_),
    .B1(_1790_),
    .B2(net194),
    .C1(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__o21a_1 _4939_ (.A1(_1694_),
    .A2(_1794_),
    .B1(_0997_),
    .X(_0187_));
 sky130_fd_sc_hd__or4_2 _4940_ (.A(_0791_),
    .B(_0907_),
    .C(_0694_),
    .D(_1211_),
    .X(_1795_));
 sky130_fd_sc_hd__nor2_1 _4941_ (.A(_0744_),
    .B(_1795_),
    .Y(_1796_));
 sky130_fd_sc_hd__nor2_8 _4942_ (.A(\core_0.execute.alu_mul_div.cbit[0] ),
    .B(\core_0.execute.alu_mul_div.cbit[1] ),
    .Y(_1797_));
 sky130_fd_sc_hd__nor2_1 _4943_ (.A(_1437_),
    .B(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__a22o_1 _4944_ (.A1(_1207_),
    .A2(_1795_),
    .B1(_1796_),
    .B2(_1798_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_4 _4945_ (.A(_1204_),
    .X(_1799_));
 sky130_fd_sc_hd__nor2_1 _4946_ (.A(_1436_),
    .B(_1437_),
    .Y(_1800_));
 sky130_fd_sc_hd__or4b_1 _4947_ (.A(_0744_),
    .B(_1209_),
    .C(_1800_),
    .D_N(_1212_),
    .X(_1801_));
 sky130_fd_sc_hd__o21ai_1 _4948_ (.A1(_1799_),
    .A2(_1212_),
    .B1(_1801_),
    .Y(_0189_));
 sky130_fd_sc_hd__clkinv_2 _4949_ (.A(\core_0.execute.alu_mul_div.cbit[3] ),
    .Y(_1802_));
 sky130_fd_sc_hd__buf_4 _4950_ (.A(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__xnor2_1 _4951_ (.A(_1803_),
    .B(_1209_),
    .Y(_1804_));
 sky130_fd_sc_hd__a22o_1 _4952_ (.A1(_1202_),
    .A2(_1795_),
    .B1(_1796_),
    .B2(_1804_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _4953_ (.A0(\core_0.de_jmp_pred ),
    .A1(\core_0.decode.i_jmp_pred_pass ),
    .S(_0913_),
    .X(_1805_));
 sky130_fd_sc_hd__clkbuf_1 _4954_ (.A(_1805_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _4955_ (.A0(\core_0.execute.sreg_data_page ),
    .A1(net104),
    .S(_0740_),
    .X(_1806_));
 sky130_fd_sc_hd__and2_1 _4956_ (.A(_1190_),
    .B(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__clkbuf_1 _4957_ (.A(_1807_),
    .X(_0192_));
 sky130_fd_sc_hd__or4_1 _4958_ (.A(net72),
    .B(_1069_),
    .C(_1070_),
    .D(_0697_),
    .X(_1808_));
 sky130_fd_sc_hd__o211a_1 _4959_ (.A1(\core_0.execute.mem_stage_pc[0] ),
    .A2(_1028_),
    .B1(_1808_),
    .C1(_0997_),
    .X(_0193_));
 sky130_fd_sc_hd__or4_1 _4960_ (.A(net79),
    .B(_1069_),
    .C(_1070_),
    .D(_0697_),
    .X(_1809_));
 sky130_fd_sc_hd__o211a_1 _4961_ (.A1(\core_0.execute.mem_stage_pc[1] ),
    .A2(_1028_),
    .B1(_1809_),
    .C1(_0997_),
    .X(_0194_));
 sky130_fd_sc_hd__or4_1 _4962_ (.A(net80),
    .B(_1069_),
    .C(_1070_),
    .D(_0697_),
    .X(_1810_));
 sky130_fd_sc_hd__o211a_1 _4963_ (.A1(\core_0.execute.mem_stage_pc[2] ),
    .A2(_1028_),
    .B1(_1810_),
    .C1(_0997_),
    .X(_0195_));
 sky130_fd_sc_hd__or4_1 _4964_ (.A(net81),
    .B(_1069_),
    .C(_1070_),
    .D(_0697_),
    .X(_1811_));
 sky130_fd_sc_hd__o211a_1 _4965_ (.A1(\core_0.execute.mem_stage_pc[3] ),
    .A2(_1028_),
    .B1(_1811_),
    .C1(_0997_),
    .X(_0196_));
 sky130_fd_sc_hd__or4_1 _4966_ (.A(net82),
    .B(_1069_),
    .C(_1070_),
    .D(_0697_),
    .X(_1812_));
 sky130_fd_sc_hd__o211a_1 _4967_ (.A1(\core_0.execute.mem_stage_pc[4] ),
    .A2(_1028_),
    .B1(_1812_),
    .C1(_0997_),
    .X(_0197_));
 sky130_fd_sc_hd__inv_2 _4968_ (.A(net83),
    .Y(_1813_));
 sky130_fd_sc_hd__buf_4 _4969_ (.A(_1027_),
    .X(_1814_));
 sky130_fd_sc_hd__nand2_1 _4970_ (.A(_1813_),
    .B(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__o211a_1 _4971_ (.A1(\core_0.execute.mem_stage_pc[5] ),
    .A2(_1028_),
    .B1(_1815_),
    .C1(_0997_),
    .X(_0198_));
 sky130_fd_sc_hd__inv_2 _4972_ (.A(net84),
    .Y(_1816_));
 sky130_fd_sc_hd__nand2_1 _4973_ (.A(_1816_),
    .B(_1814_),
    .Y(_1817_));
 sky130_fd_sc_hd__buf_4 _4974_ (.A(_1314_),
    .X(_1818_));
 sky130_fd_sc_hd__o211a_1 _4975_ (.A1(\core_0.execute.mem_stage_pc[6] ),
    .A2(_1028_),
    .B1(_1817_),
    .C1(_1818_),
    .X(_0199_));
 sky130_fd_sc_hd__inv_2 _4976_ (.A(net85),
    .Y(_1819_));
 sky130_fd_sc_hd__nand2_1 _4977_ (.A(_1819_),
    .B(_1814_),
    .Y(_1820_));
 sky130_fd_sc_hd__o211a_1 _4978_ (.A1(\core_0.execute.mem_stage_pc[7] ),
    .A2(_1028_),
    .B1(_1820_),
    .C1(_1818_),
    .X(_0200_));
 sky130_fd_sc_hd__or4_1 _4979_ (.A(net86),
    .B(_1069_),
    .C(_1070_),
    .D(_0697_),
    .X(_1821_));
 sky130_fd_sc_hd__o211a_1 _4980_ (.A1(\core_0.execute.mem_stage_pc[8] ),
    .A2(_1028_),
    .B1(_1821_),
    .C1(_1818_),
    .X(_0201_));
 sky130_fd_sc_hd__or4_1 _4981_ (.A(net87),
    .B(_1069_),
    .C(_1070_),
    .D(_0697_),
    .X(_1822_));
 sky130_fd_sc_hd__o211a_1 _4982_ (.A1(\core_0.execute.mem_stage_pc[9] ),
    .A2(_1814_),
    .B1(_1822_),
    .C1(_1818_),
    .X(_0202_));
 sky130_fd_sc_hd__inv_2 _4983_ (.A(net73),
    .Y(_1823_));
 sky130_fd_sc_hd__nand2_1 _4984_ (.A(_1823_),
    .B(_1027_),
    .Y(_1824_));
 sky130_fd_sc_hd__o211a_1 _4985_ (.A1(\core_0.execute.mem_stage_pc[10] ),
    .A2(_1814_),
    .B1(_1824_),
    .C1(_1818_),
    .X(_0203_));
 sky130_fd_sc_hd__inv_2 _4986_ (.A(net74),
    .Y(_1825_));
 sky130_fd_sc_hd__nand2_1 _4987_ (.A(_1825_),
    .B(_1027_),
    .Y(_1826_));
 sky130_fd_sc_hd__o211a_1 _4988_ (.A1(\core_0.execute.mem_stage_pc[11] ),
    .A2(_1814_),
    .B1(_1826_),
    .C1(_1818_),
    .X(_0204_));
 sky130_fd_sc_hd__or4_1 _4989_ (.A(net75),
    .B(_1069_),
    .C(_1070_),
    .D(_0697_),
    .X(_1827_));
 sky130_fd_sc_hd__o211a_1 _4990_ (.A1(\core_0.execute.mem_stage_pc[12] ),
    .A2(_1814_),
    .B1(_1827_),
    .C1(_1818_),
    .X(_0205_));
 sky130_fd_sc_hd__inv_2 _4991_ (.A(net76),
    .Y(_1828_));
 sky130_fd_sc_hd__nand2_1 _4992_ (.A(_1828_),
    .B(_1027_),
    .Y(_1829_));
 sky130_fd_sc_hd__o211a_1 _4993_ (.A1(\core_0.execute.mem_stage_pc[13] ),
    .A2(_1814_),
    .B1(_1829_),
    .C1(_1818_),
    .X(_0206_));
 sky130_fd_sc_hd__inv_2 _4994_ (.A(net77),
    .Y(_1830_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(_1830_),
    .B(_1027_),
    .Y(_1831_));
 sky130_fd_sc_hd__o211a_1 _4996_ (.A1(\core_0.execute.mem_stage_pc[14] ),
    .A2(_1814_),
    .B1(_1831_),
    .C1(_1818_),
    .X(_0207_));
 sky130_fd_sc_hd__or4_1 _4997_ (.A(net78),
    .B(_1069_),
    .C(_1070_),
    .D(_0697_),
    .X(_1832_));
 sky130_fd_sc_hd__o211a_1 _4998_ (.A1(\core_0.execute.mem_stage_pc[15] ),
    .A2(_1814_),
    .B1(_1832_),
    .C1(_1818_),
    .X(_0208_));
 sky130_fd_sc_hd__nor2_1 _4999_ (.A(_1128_),
    .B(_0689_),
    .Y(_0209_));
 sky130_fd_sc_hd__nor2_1 _5000_ (.A(_1128_),
    .B(_0687_),
    .Y(_0210_));
 sky130_fd_sc_hd__nor2_1 _5001_ (.A(_1128_),
    .B(_0676_),
    .Y(_0211_));
 sky130_fd_sc_hd__nor2_1 _5002_ (.A(_1128_),
    .B(_0678_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor2_1 _5003_ (.A(_1128_),
    .B(_0682_),
    .Y(_0213_));
 sky130_fd_sc_hd__nor2_1 _5004_ (.A(_1128_),
    .B(_0685_),
    .Y(_0214_));
 sky130_fd_sc_hd__nor2_1 _5005_ (.A(_1157_),
    .B(_0681_),
    .Y(_0215_));
 sky130_fd_sc_hd__nor2_1 _5006_ (.A(_1157_),
    .B(_0677_),
    .Y(_0216_));
 sky130_fd_sc_hd__and3_1 _5007_ (.A(\core_0.execute.trap_flag ),
    .B(_0996_),
    .C(_1071_),
    .X(_1833_));
 sky130_fd_sc_hd__clkbuf_1 _5008_ (.A(_1833_),
    .X(_0217_));
 sky130_fd_sc_hd__and3_2 _5009_ (.A(\core_0.dec_sys ),
    .B(_0995_),
    .C(_1071_),
    .X(_1834_));
 sky130_fd_sc_hd__clkbuf_1 _5010_ (.A(_1834_),
    .X(_0218_));
 sky130_fd_sc_hd__nand2_4 _5011_ (.A(_0665_),
    .B(_1027_),
    .Y(_1835_));
 sky130_fd_sc_hd__clkbuf_8 _5012_ (.A(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__mux2_1 _5013_ (.A0(\core_0.dec_mem_we ),
    .A1(net159),
    .S(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__clkbuf_1 _5014_ (.A(_1837_),
    .X(_0219_));
 sky130_fd_sc_hd__or4_4 _5015_ (.A(_1636_),
    .B(_1640_),
    .C(_1641_),
    .D(_1642_),
    .X(_1838_));
 sky130_fd_sc_hd__or2_4 _5016_ (.A(_1323_),
    .B(_1325_),
    .X(_1839_));
 sky130_fd_sc_hd__nor2_2 _5017_ (.A(_1332_),
    .B(_1609_),
    .Y(_1840_));
 sky130_fd_sc_hd__o22a_4 _5018_ (.A1(net93),
    .A2(_1572_),
    .B1(_1604_),
    .B2(_1608_),
    .X(_1841_));
 sky130_fd_sc_hd__nor2_1 _5019_ (.A(_1331_),
    .B(_1841_),
    .Y(_1842_));
 sky130_fd_sc_hd__nor2_2 _5020_ (.A(_1840_),
    .B(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__or3_1 _5021_ (.A(_1334_),
    .B(_1601_),
    .C(_1843_),
    .X(_1844_));
 sky130_fd_sc_hd__a21o_1 _5022_ (.A1(_1077_),
    .A2(net182),
    .B1(_1333_),
    .X(_1845_));
 sky130_fd_sc_hd__nor2_1 _5023_ (.A(_1845_),
    .B(_1601_),
    .Y(_1846_));
 sky130_fd_sc_hd__nor2_2 _5024_ (.A(_1334_),
    .B(_1757_),
    .Y(_1847_));
 sky130_fd_sc_hd__nor2_2 _5025_ (.A(_1846_),
    .B(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__o21a_1 _5026_ (.A1(_1338_),
    .A2(_1588_),
    .B1(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__or3_1 _5027_ (.A(_1338_),
    .B(_1588_),
    .C(_1848_),
    .X(_1850_));
 sky130_fd_sc_hd__and2b_1 _5028_ (.A_N(_1849_),
    .B(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__nor2_2 _5029_ (.A(_1338_),
    .B(_1756_),
    .Y(_1852_));
 sky130_fd_sc_hd__nand2_1 _5030_ (.A(_1338_),
    .B(_1756_),
    .Y(_1853_));
 sky130_fd_sc_hd__and2b_1 _5031_ (.A_N(_1852_),
    .B(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__nor2_1 _5032_ (.A(_1594_),
    .B(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__o21a_1 _5033_ (.A1(_1342_),
    .A2(_1594_),
    .B1(_1854_),
    .X(_1856_));
 sky130_fd_sc_hd__a21oi_2 _5034_ (.A1(_1493_),
    .A2(_1855_),
    .B1(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__or2_1 _5035_ (.A(_1482_),
    .B(_1549_),
    .X(_1858_));
 sky130_fd_sc_hd__nand2_1 _5036_ (.A(_1482_),
    .B(_1549_),
    .Y(_1859_));
 sky130_fd_sc_hd__and2_1 _5037_ (.A(_1858_),
    .B(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__o21a_1 _5038_ (.A1(_1392_),
    .A2(_1579_),
    .B1(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__o22ai_4 _5039_ (.A1(net102),
    .A2(_1572_),
    .B1(_1573_),
    .B2(_1578_),
    .Y(_1862_));
 sky130_fd_sc_hd__and3b_1 _5040_ (.A_N(_1860_),
    .B(_1391_),
    .C(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__nor2_1 _5041_ (.A(_1861_),
    .B(_1863_),
    .Y(_1864_));
 sky130_fd_sc_hd__nor2_1 _5042_ (.A(_1353_),
    .B(_1745_),
    .Y(_1865_));
 sky130_fd_sc_hd__nand2_1 _5043_ (.A(_1353_),
    .B(_1745_),
    .Y(_1866_));
 sky130_fd_sc_hd__nand2b_1 _5044_ (.A_N(_1865_),
    .B(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__a21oi_1 _5045_ (.A1(_1357_),
    .A2(_1746_),
    .B1(_1867_),
    .Y(_1868_));
 sky130_fd_sc_hd__and3_1 _5046_ (.A(_1357_),
    .B(_1746_),
    .C(_1867_),
    .X(_1869_));
 sky130_fd_sc_hd__nor2_1 _5047_ (.A(_1868_),
    .B(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__and2_1 _5048_ (.A(_1357_),
    .B(_1654_),
    .X(_1871_));
 sky130_fd_sc_hd__nor2_1 _5049_ (.A(_1357_),
    .B(_1654_),
    .Y(_1872_));
 sky130_fd_sc_hd__nor2_2 _5050_ (.A(_1871_),
    .B(_1872_),
    .Y(_1873_));
 sky130_fd_sc_hd__nor2_1 _5051_ (.A(_1661_),
    .B(_1873_),
    .Y(_1874_));
 sky130_fd_sc_hd__o21a_1 _5052_ (.A1(_1362_),
    .A2(_1661_),
    .B1(_1873_),
    .X(_1875_));
 sky130_fd_sc_hd__a21oi_1 _5053_ (.A1(_1709_),
    .A2(_1874_),
    .B1(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__xnor2_4 _5054_ (.A(_1362_),
    .B(_1743_),
    .Y(_1877_));
 sky130_fd_sc_hd__a21oi_1 _5055_ (.A1(_1701_),
    .A2(_1677_),
    .B1(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__nand3_1 _5056_ (.A(_1701_),
    .B(_1677_),
    .C(_1877_),
    .Y(_1879_));
 sky130_fd_sc_hd__and2b_1 _5057_ (.A_N(_1878_),
    .B(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__nand2_1 _5058_ (.A(_1698_),
    .B(_1633_),
    .Y(_1881_));
 sky130_fd_sc_hd__o22a_1 _5059_ (.A1(_1419_),
    .A2(_1420_),
    .B1(_1766_),
    .B2(_1763_),
    .X(_1882_));
 sky130_fd_sc_hd__and2_1 _5060_ (.A(_1766_),
    .B(_1763_),
    .X(_1883_));
 sky130_fd_sc_hd__o21ai_1 _5061_ (.A1(_1882_),
    .A2(_1883_),
    .B1(_1624_),
    .Y(_1884_));
 sky130_fd_sc_hd__or3_1 _5062_ (.A(_1624_),
    .B(_1882_),
    .C(_1883_),
    .X(_1885_));
 sky130_fd_sc_hd__a21bo_2 _5063_ (.A1(_1738_),
    .A2(_1884_),
    .B1_N(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__nor2_1 _5064_ (.A(_1698_),
    .B(_1633_),
    .Y(_1887_));
 sky130_fd_sc_hd__nor2_1 _5065_ (.A(_1370_),
    .B(_1670_),
    .Y(_1888_));
 sky130_fd_sc_hd__nand2_1 _5066_ (.A(_1370_),
    .B(_1670_),
    .Y(_1889_));
 sky130_fd_sc_hd__nor2b_1 _5067_ (.A(_1888_),
    .B_N(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__a211o_1 _5068_ (.A1(_1881_),
    .A2(_1886_),
    .B1(_1887_),
    .C1(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__nor2_1 _5069_ (.A(_1365_),
    .B(_1676_),
    .Y(_1892_));
 sky130_fd_sc_hd__nand2_1 _5070_ (.A(_1365_),
    .B(_1677_),
    .Y(_1893_));
 sky130_fd_sc_hd__and2b_1 _5071_ (.A_N(_1892_),
    .B(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__clkbuf_4 _5072_ (.A(_1894_),
    .X(_1895_));
 sky130_fd_sc_hd__nand2_1 _5073_ (.A(_1703_),
    .B(_1670_),
    .Y(_1896_));
 sky130_fd_sc_hd__xor2_1 _5074_ (.A(_1895_),
    .B(_1896_),
    .X(_1897_));
 sky130_fd_sc_hd__a31o_1 _5075_ (.A1(_1879_),
    .A2(_1895_),
    .A3(_1896_),
    .B1(_1878_),
    .X(_1898_));
 sky130_fd_sc_hd__a31o_1 _5076_ (.A1(_1880_),
    .A2(_1891_),
    .A3(_1897_),
    .B1(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__o21ba_1 _5077_ (.A1(_1868_),
    .A2(_1875_),
    .B1_N(_1869_),
    .X(_1900_));
 sky130_fd_sc_hd__a31o_1 _5078_ (.A1(_1870_),
    .A2(_1876_),
    .A3(_1899_),
    .B1(_1900_),
    .X(_1901_));
 sky130_fd_sc_hd__a21o_2 _5079_ (.A1(_1077_),
    .A2(net191),
    .B1(_1352_),
    .X(_1902_));
 sky130_fd_sc_hd__nor2_2 _5080_ (.A(_1392_),
    .B(_1862_),
    .Y(_1903_));
 sky130_fd_sc_hd__or2_1 _5081_ (.A(_1391_),
    .B(_1579_),
    .X(_1904_));
 sky130_fd_sc_hd__nor2b_2 _5082_ (.A(_1903_),
    .B_N(_1904_),
    .Y(_1905_));
 sky130_fd_sc_hd__nor2_1 _5083_ (.A(_1571_),
    .B(_1905_),
    .Y(_1906_));
 sky130_fd_sc_hd__o21a_1 _5084_ (.A1(_1353_),
    .A2(_1571_),
    .B1(_1905_),
    .X(_1907_));
 sky130_fd_sc_hd__a21oi_1 _5085_ (.A1(_1902_),
    .A2(_1906_),
    .B1(_1907_),
    .Y(_1908_));
 sky130_fd_sc_hd__inv_2 _5086_ (.A(_1863_),
    .Y(_1909_));
 sky130_fd_sc_hd__a21o_1 _5087_ (.A1(_1909_),
    .A2(_1907_),
    .B1(_1861_),
    .X(_1910_));
 sky130_fd_sc_hd__a31o_1 _5088_ (.A1(_1864_),
    .A2(_1901_),
    .A3(_1908_),
    .B1(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__or2_1 _5089_ (.A(_1493_),
    .B(_1594_),
    .X(_1912_));
 sky130_fd_sc_hd__inv_2 _5090_ (.A(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__o22ai_4 _5091_ (.A1(net90),
    .A2(_1572_),
    .B1(_1590_),
    .B2(_1593_),
    .Y(_1914_));
 sky130_fd_sc_hd__nor2_1 _5092_ (.A(_1342_),
    .B(_1914_),
    .Y(_1915_));
 sky130_fd_sc_hd__nor2_2 _5093_ (.A(_1913_),
    .B(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hd__o21a_1 _5094_ (.A1(_1345_),
    .A2(_1558_),
    .B1(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__or3_1 _5095_ (.A(_1345_),
    .B(_1558_),
    .C(_1916_),
    .X(_1918_));
 sky130_fd_sc_hd__or2b_1 _5096_ (.A(_1917_),
    .B_N(_1918_),
    .X(_1919_));
 sky130_fd_sc_hd__clkinv_2 _5097_ (.A(_1557_),
    .Y(_1920_));
 sky130_fd_sc_hd__nor2_2 _5098_ (.A(_1345_),
    .B(_1920_),
    .Y(_1921_));
 sky130_fd_sc_hd__or2_1 _5099_ (.A(_1344_),
    .B(_1558_),
    .X(_1922_));
 sky130_fd_sc_hd__and2b_1 _5100_ (.A_N(_1921_),
    .B(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__nor2_1 _5101_ (.A(_1550_),
    .B(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__o21a_1 _5102_ (.A1(_1350_),
    .A2(_1550_),
    .B1(_1923_),
    .X(_1925_));
 sky130_fd_sc_hd__a21o_1 _5103_ (.A1(_1482_),
    .A2(_1924_),
    .B1(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__nor2_1 _5104_ (.A(_1919_),
    .B(_1926_),
    .Y(_1927_));
 sky130_fd_sc_hd__or2_1 _5105_ (.A(_1917_),
    .B(_1925_),
    .X(_1928_));
 sky130_fd_sc_hd__a22o_1 _5106_ (.A1(_1911_),
    .A2(_1927_),
    .B1(_1928_),
    .B2(_1918_),
    .X(_1929_));
 sky130_fd_sc_hd__o21a_1 _5107_ (.A1(_1849_),
    .A2(_1856_),
    .B1(_1850_),
    .X(_1930_));
 sky130_fd_sc_hd__a31o_1 _5108_ (.A1(_1851_),
    .A2(_1857_),
    .A3(_1929_),
    .B1(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__nand2_1 _5109_ (.A(_1326_),
    .B(_1541_),
    .Y(_1932_));
 sky130_fd_sc_hd__or2_1 _5110_ (.A(_1326_),
    .B(_1541_),
    .X(_1933_));
 sky130_fd_sc_hd__and2_1 _5111_ (.A(_1932_),
    .B(_1933_),
    .X(_1934_));
 sky130_fd_sc_hd__o21a_1 _5112_ (.A1(_1332_),
    .A2(_1841_),
    .B1(_1934_),
    .X(_1935_));
 sky130_fd_sc_hd__o21a_1 _5113_ (.A1(_1334_),
    .A2(_1601_),
    .B1(_1843_),
    .X(_1936_));
 sky130_fd_sc_hd__a211oi_1 _5114_ (.A1(_1844_),
    .A2(_1931_),
    .B1(_1935_),
    .C1(_1936_),
    .Y(_1937_));
 sky130_fd_sc_hd__and3b_1 _5115_ (.A_N(_1934_),
    .B(_1331_),
    .C(_1609_),
    .X(_1938_));
 sky130_fd_sc_hd__a211o_1 _5116_ (.A1(_1839_),
    .A2(_1541_),
    .B1(_1937_),
    .C1(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__nor2_1 _5117_ (.A(_1326_),
    .B(_1541_),
    .Y(_1940_));
 sky130_fd_sc_hd__or2_1 _5118_ (.A(_1915_),
    .B(_1921_),
    .X(_1941_));
 sky130_fd_sc_hd__nand2_1 _5119_ (.A(_1374_),
    .B(_1633_),
    .Y(_1942_));
 sky130_fd_sc_hd__nand2_1 _5120_ (.A(_1738_),
    .B(_1624_),
    .Y(_1943_));
 sky130_fd_sc_hd__a21o_1 _5121_ (.A1(_1736_),
    .A2(_1763_),
    .B1(_1767_),
    .X(_1944_));
 sky130_fd_sc_hd__nor2_1 _5122_ (.A(_1374_),
    .B(_1632_),
    .Y(_1945_));
 sky130_fd_sc_hd__nor2_1 _5123_ (.A(_1738_),
    .B(_1624_),
    .Y(_1946_));
 sky130_fd_sc_hd__a211o_1 _5124_ (.A1(_1943_),
    .A2(_1944_),
    .B1(_1945_),
    .C1(_1946_),
    .X(_1947_));
 sky130_fd_sc_hd__a31o_1 _5125_ (.A1(_1889_),
    .A2(_1942_),
    .A3(_1947_),
    .B1(_1888_),
    .X(_1948_));
 sky130_fd_sc_hd__and2b_1 _5126_ (.A_N(_1865_),
    .B(_1866_),
    .X(_1949_));
 sky130_fd_sc_hd__and2_1 _5127_ (.A(_1949_),
    .B(_1873_),
    .X(_1950_));
 sky130_fd_sc_hd__and4b_1 _5128_ (.A_N(_1877_),
    .B(_1895_),
    .C(_1948_),
    .D(_1950_),
    .X(_1951_));
 sky130_fd_sc_hd__nor2_1 _5129_ (.A(_1362_),
    .B(_1743_),
    .Y(_1952_));
 sky130_fd_sc_hd__nand2_1 _5130_ (.A(_1362_),
    .B(_1743_),
    .Y(_1953_));
 sky130_fd_sc_hd__o21a_1 _5131_ (.A1(_1952_),
    .A2(_1892_),
    .B1(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__or2_1 _5132_ (.A(_1357_),
    .B(_1654_),
    .X(_1955_));
 sky130_fd_sc_hd__o211a_1 _5133_ (.A1(_1871_),
    .A2(_1954_),
    .B1(_1955_),
    .C1(_1866_),
    .X(_1956_));
 sky130_fd_sc_hd__o31a_2 _5134_ (.A1(_1865_),
    .A2(_1951_),
    .A3(_1956_),
    .B1(_1905_),
    .X(_1957_));
 sky130_fd_sc_hd__inv_2 _5135_ (.A(_1859_),
    .Y(_1958_));
 sky130_fd_sc_hd__or2_1 _5136_ (.A(_1958_),
    .B(_1903_),
    .X(_1959_));
 sky130_fd_sc_hd__o211a_1 _5137_ (.A1(_1957_),
    .A2(_1959_),
    .B1(_1858_),
    .C1(_1923_),
    .X(_1960_));
 sky130_fd_sc_hd__o211a_1 _5138_ (.A1(_1941_),
    .A2(_1960_),
    .B1(_1854_),
    .C1(_1912_),
    .X(_1961_));
 sky130_fd_sc_hd__nand2_1 _5139_ (.A(_1334_),
    .B(_1757_),
    .Y(_1962_));
 sky130_fd_sc_hd__o311a_1 _5140_ (.A1(_1847_),
    .A2(_1852_),
    .A3(_1961_),
    .B1(_1962_),
    .C1(_1843_),
    .X(_1963_));
 sky130_fd_sc_hd__o311a_1 _5141_ (.A1(_1940_),
    .A2(_1840_),
    .A3(_1963_),
    .B1(_1932_),
    .C1(_0962_),
    .X(_1964_));
 sky130_fd_sc_hd__buf_2 _5142_ (.A(_1702_),
    .X(_1965_));
 sky130_fd_sc_hd__or2_2 _5143_ (.A(_1965_),
    .B(_1700_),
    .X(_1966_));
 sky130_fd_sc_hd__xnor2_4 _5144_ (.A(_1371_),
    .B(_1966_),
    .Y(_1967_));
 sky130_fd_sc_hd__a211o_1 _5145_ (.A1(_1965_),
    .A2(_1746_),
    .B1(_1719_),
    .C1(_1721_),
    .X(_1968_));
 sky130_fd_sc_hd__a211o_1 _5146_ (.A1(_1965_),
    .A2(_1743_),
    .B1(_1719_),
    .C1(_1721_),
    .X(_1969_));
 sky130_fd_sc_hd__mux2_1 _5147_ (.A0(_1968_),
    .A1(_1969_),
    .S(_1764_),
    .X(_1970_));
 sky130_fd_sc_hd__a211o_1 _5148_ (.A1(_1965_),
    .A2(_1745_),
    .B1(_1719_),
    .C1(_1721_),
    .X(_1971_));
 sky130_fd_sc_hd__a211o_1 _5149_ (.A1(_1965_),
    .A2(_1862_),
    .B1(_1718_),
    .C1(_1720_),
    .X(_1972_));
 sky130_fd_sc_hd__mux2_1 _5150_ (.A0(_1971_),
    .A1(_1972_),
    .S(_1422_),
    .X(_1973_));
 sky130_fd_sc_hd__nand2_2 _5151_ (.A(\core_0.decode.oc_alu_mode[12] ),
    .B(_1729_),
    .Y(_1974_));
 sky130_fd_sc_hd__xnor2_4 _5152_ (.A(_1738_),
    .B(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__mux2_1 _5153_ (.A0(_1970_),
    .A1(_1973_),
    .S(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__a211o_1 _5154_ (.A1(_1965_),
    .A2(_1677_),
    .B1(_1719_),
    .C1(_1721_),
    .X(_1977_));
 sky130_fd_sc_hd__a211o_1 _5155_ (.A1(_1965_),
    .A2(_1670_),
    .B1(_1719_),
    .C1(_1721_),
    .X(_1978_));
 sky130_fd_sc_hd__a211o_1 _5156_ (.A1(_1965_),
    .A2(_1633_),
    .B1(_1718_),
    .C1(_1720_),
    .X(_1979_));
 sky130_fd_sc_hd__a211o_1 _5157_ (.A1(_1965_),
    .A2(_1624_),
    .B1(_1719_),
    .C1(_1721_),
    .X(_1980_));
 sky130_fd_sc_hd__xnor2_2 _5158_ (.A(_1725_),
    .B(_1974_),
    .Y(_1981_));
 sky130_fd_sc_hd__mux4_1 _5159_ (.A0(_1977_),
    .A1(_1978_),
    .A2(_1979_),
    .A3(_1980_),
    .S0(_1764_),
    .S1(_1981_),
    .X(_1982_));
 sky130_fd_sc_hd__nor2_2 _5160_ (.A(_1724_),
    .B(_1764_),
    .Y(_1983_));
 sky130_fd_sc_hd__nor2_2 _5161_ (.A(_1965_),
    .B(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__xnor2_1 _5162_ (.A(_1374_),
    .B(_1984_),
    .Y(_1985_));
 sky130_fd_sc_hd__mux2_1 _5163_ (.A0(_1976_),
    .A1(_1982_),
    .S(_1985_),
    .X(_1986_));
 sky130_fd_sc_hd__nor2_1 _5164_ (.A(_1967_),
    .B(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__xnor2_4 _5165_ (.A(_1749_),
    .B(_1984_),
    .Y(_1988_));
 sky130_fd_sc_hd__o21a_1 _5166_ (.A1(_0984_),
    .A2(_1594_),
    .B1(_1722_),
    .X(_1989_));
 sky130_fd_sc_hd__o21a_1 _5167_ (.A1(_0984_),
    .A2(_1588_),
    .B1(_1722_),
    .X(_1990_));
 sky130_fd_sc_hd__mux2_1 _5168_ (.A0(_1989_),
    .A1(_1990_),
    .S(_1423_),
    .X(_1991_));
 sky130_fd_sc_hd__o21a_1 _5169_ (.A1(_0984_),
    .A2(_1558_),
    .B1(_1722_),
    .X(_1992_));
 sky130_fd_sc_hd__nor4_4 _5170_ (.A(_1713_),
    .B(_1714_),
    .C(_1734_),
    .D(_1717_),
    .Y(_1993_));
 sky130_fd_sc_hd__nand2_1 _5171_ (.A(_0984_),
    .B(_1541_),
    .Y(_1994_));
 sky130_fd_sc_hd__o211ai_2 _5172_ (.A1(_0984_),
    .A2(_1550_),
    .B1(_1993_),
    .C1(_1994_),
    .Y(_1995_));
 sky130_fd_sc_hd__nor2_1 _5173_ (.A(_1422_),
    .B(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__a21o_1 _5174_ (.A1(_1423_),
    .A2(_1992_),
    .B1(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__clkbuf_4 _5175_ (.A(_1981_),
    .X(_1998_));
 sky130_fd_sc_hd__mux2_1 _5176_ (.A0(_1991_),
    .A1(_1997_),
    .S(_1998_),
    .X(_1999_));
 sky130_fd_sc_hd__o21a_1 _5177_ (.A1(_0984_),
    .A2(_1841_),
    .B1(_1722_),
    .X(_2000_));
 sky130_fd_sc_hd__o21a_1 _5178_ (.A1(_0984_),
    .A2(_1601_),
    .B1(_1722_),
    .X(_2001_));
 sky130_fd_sc_hd__buf_4 _5179_ (.A(_1764_),
    .X(_2002_));
 sky130_fd_sc_hd__mux2_1 _5180_ (.A0(_2000_),
    .A1(_2001_),
    .S(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__nand2_1 _5181_ (.A(_1542_),
    .B(_1993_),
    .Y(_2004_));
 sky130_fd_sc_hd__nor2_1 _5182_ (.A(_2004_),
    .B(_1998_),
    .Y(_2005_));
 sky130_fd_sc_hd__buf_2 _5183_ (.A(_1985_),
    .X(_2006_));
 sky130_fd_sc_hd__a221o_1 _5184_ (.A1(_1998_),
    .A2(_2003_),
    .B1(_2005_),
    .B2(_2002_),
    .C1(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__o211a_1 _5185_ (.A1(_1988_),
    .A2(_1999_),
    .B1(_2007_),
    .C1(_1967_),
    .X(_2008_));
 sky130_fd_sc_hd__nand2_1 _5186_ (.A(_1371_),
    .B(_1700_),
    .Y(_2009_));
 sky130_fd_sc_hd__or3_1 _5187_ (.A(_1708_),
    .B(_1719_),
    .C(_1721_),
    .X(_2010_));
 sky130_fd_sc_hd__o21ai_1 _5188_ (.A1(_2009_),
    .A2(_2010_),
    .B1(_1705_),
    .Y(_2011_));
 sky130_fd_sc_hd__o211a_1 _5189_ (.A1(_1362_),
    .A2(_1714_),
    .B1(_2011_),
    .C1(\core_0.decode.oc_alu_mode[13] ),
    .X(_2012_));
 sky130_fd_sc_hd__o31a_1 _5190_ (.A1(_1705_),
    .A2(_1987_),
    .A3(_2008_),
    .B1(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__a211oi_4 _5191_ (.A1(_0978_),
    .A2(_1939_),
    .B1(_1964_),
    .C1(_2013_),
    .Y(_2014_));
 sky130_fd_sc_hd__nand2_1 _5192_ (.A(_1326_),
    .B(_2014_),
    .Y(_2015_));
 sky130_fd_sc_hd__xor2_1 _5193_ (.A(_1838_),
    .B(_2015_),
    .X(_2016_));
 sky130_fd_sc_hd__mux2_1 _5194_ (.A0(_2016_),
    .A1(\core_0.ew_addr_high[0] ),
    .S(_1836_),
    .X(_2017_));
 sky130_fd_sc_hd__clkbuf_1 _5195_ (.A(_2017_),
    .X(_0220_));
 sky130_fd_sc_hd__nand4_4 _5196_ (.A(_1614_),
    .B(_1618_),
    .C(_1619_),
    .D(_1620_),
    .Y(_2018_));
 sky130_fd_sc_hd__or2_1 _5197_ (.A(_1838_),
    .B(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__nand2_1 _5198_ (.A(_1838_),
    .B(_2018_),
    .Y(_2020_));
 sky130_fd_sc_hd__nand2_2 _5199_ (.A(_2019_),
    .B(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__o21a_1 _5200_ (.A1(_1839_),
    .A2(_1838_),
    .B1(_2014_),
    .X(_2022_));
 sky130_fd_sc_hd__xnor2_4 _5201_ (.A(_2021_),
    .B(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__mux2_1 _5202_ (.A0(_2023_),
    .A1(net132),
    .S(_1836_),
    .X(_2024_));
 sky130_fd_sc_hd__clkbuf_1 _5203_ (.A(_2024_),
    .X(_0221_));
 sky130_fd_sc_hd__nand2_2 _5204_ (.A(_1839_),
    .B(_2014_),
    .Y(_2025_));
 sky130_fd_sc_hd__a22o_2 _5205_ (.A1(_2014_),
    .A2(_2019_),
    .B1(_2020_),
    .B2(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__nor2_4 _5206_ (.A(_1630_),
    .B(_1626_),
    .Y(_2027_));
 sky130_fd_sc_hd__xor2_4 _5207_ (.A(_2026_),
    .B(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__mux2_1 _5208_ (.A0(_2028_),
    .A1(net133),
    .S(_1836_),
    .X(_2029_));
 sky130_fd_sc_hd__clkbuf_1 _5209_ (.A(_2029_),
    .X(_0222_));
 sky130_fd_sc_hd__and2b_1 _5210_ (.A_N(_2019_),
    .B(_2027_),
    .X(_2030_));
 sky130_fd_sc_hd__or2b_1 _5211_ (.A(_2025_),
    .B_N(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__or3_1 _5212_ (.A(_2014_),
    .B(_2020_),
    .C(_2027_),
    .X(_2032_));
 sky130_fd_sc_hd__nor2_2 _5213_ (.A(_1667_),
    .B(_1665_),
    .Y(_2033_));
 sky130_fd_sc_hd__a21oi_1 _5214_ (.A1(_2031_),
    .A2(_2032_),
    .B1(_2033_),
    .Y(_2034_));
 sky130_fd_sc_hd__and3_1 _5215_ (.A(_2031_),
    .B(_2032_),
    .C(_2033_),
    .X(_2035_));
 sky130_fd_sc_hd__nor2_1 _5216_ (.A(_2034_),
    .B(_2035_),
    .Y(_2036_));
 sky130_fd_sc_hd__mux2_1 _5217_ (.A0(_2036_),
    .A1(net134),
    .S(_1836_),
    .X(_2037_));
 sky130_fd_sc_hd__clkbuf_1 _5218_ (.A(_2037_),
    .X(_0223_));
 sky130_fd_sc_hd__or2_1 _5219_ (.A(_2032_),
    .B(_2033_),
    .X(_2038_));
 sky130_fd_sc_hd__a21o_1 _5220_ (.A1(\core_0.execute.rf.reg_outputs[1][4] ),
    .A2(_1526_),
    .B1(_1674_),
    .X(_2039_));
 sky130_fd_sc_hd__nand4_1 _5221_ (.A(_1839_),
    .B(_2014_),
    .C(_2030_),
    .D(_2033_),
    .Y(_2040_));
 sky130_fd_sc_hd__and2b_1 _5222_ (.A_N(_2039_),
    .B(_2040_),
    .X(_2041_));
 sky130_fd_sc_hd__a21boi_1 _5223_ (.A1(_2038_),
    .A2(_2040_),
    .B1_N(_2039_),
    .Y(_2042_));
 sky130_fd_sc_hd__a21oi_1 _5224_ (.A1(_2038_),
    .A2(_2041_),
    .B1(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__buf_6 _5225_ (.A(_1835_),
    .X(_2044_));
 sky130_fd_sc_hd__mux2_1 _5226_ (.A0(_2043_),
    .A1(net135),
    .S(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__clkbuf_1 _5227_ (.A(_2045_),
    .X(_0224_));
 sky130_fd_sc_hd__a21o_1 _5228_ (.A1(\core_0.execute.rf.reg_outputs[1][5] ),
    .A2(_1526_),
    .B1(_1659_),
    .X(_2046_));
 sky130_fd_sc_hd__a21o_1 _5229_ (.A1(_2038_),
    .A2(_2039_),
    .B1(_2041_),
    .X(_2047_));
 sky130_fd_sc_hd__xnor2_1 _5230_ (.A(_2046_),
    .B(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__mux2_1 _5231_ (.A0(_2048_),
    .A1(net136),
    .S(_2044_),
    .X(_2049_));
 sky130_fd_sc_hd__clkbuf_1 _5232_ (.A(_2049_),
    .X(_0225_));
 sky130_fd_sc_hd__a21o_1 _5233_ (.A1(\core_0.execute.rf.reg_outputs[1][6] ),
    .A2(_1526_),
    .B1(_1649_),
    .X(_2050_));
 sky130_fd_sc_hd__xor2_1 _5234_ (.A(_2025_),
    .B(_2046_),
    .X(_2051_));
 sky130_fd_sc_hd__a211oi_1 _5235_ (.A1(_2038_),
    .A2(_2039_),
    .B1(_2041_),
    .C1(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hd__xor2_1 _5236_ (.A(_2050_),
    .B(_2052_),
    .X(_2053_));
 sky130_fd_sc_hd__mux2_1 _5237_ (.A0(_2053_),
    .A1(net137),
    .S(_2044_),
    .X(_2054_));
 sky130_fd_sc_hd__clkbuf_1 _5238_ (.A(_2054_),
    .X(_0226_));
 sky130_fd_sc_hd__a21o_1 _5239_ (.A1(\core_0.execute.rf.reg_outputs[1][7] ),
    .A2(_1526_),
    .B1(_1569_),
    .X(_2055_));
 sky130_fd_sc_hd__xor2_1 _5240_ (.A(_2025_),
    .B(_2050_),
    .X(_2056_));
 sky130_fd_sc_hd__a2111o_1 _5241_ (.A1(_2038_),
    .A2(_2039_),
    .B1(_2041_),
    .C1(_2051_),
    .D1(_2056_),
    .X(_2057_));
 sky130_fd_sc_hd__xnor2_1 _5242_ (.A(_2055_),
    .B(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__mux2_1 _5243_ (.A0(_2058_),
    .A1(net138),
    .S(_2044_),
    .X(_2059_));
 sky130_fd_sc_hd__clkbuf_1 _5244_ (.A(_2059_),
    .X(_0227_));
 sky130_fd_sc_hd__and2_1 _5245_ (.A(_0665_),
    .B(_1071_),
    .X(_2060_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _5246_ (.A(_2060_),
    .X(_0228_));
 sky130_fd_sc_hd__and2b_1 _5247_ (.A_N(net187),
    .B(net186),
    .X(_2061_));
 sky130_fd_sc_hd__and4b_1 _5248_ (.A_N(net192),
    .B(_1030_),
    .C(_1031_),
    .D(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__a31o_1 _5249_ (.A1(net185),
    .A2(_1159_),
    .A3(_2062_),
    .B1(\core_0.dec_sreg_jal_over ),
    .X(_2063_));
 sky130_fd_sc_hd__and4b_1 _5250_ (.A_N(net192),
    .B(_1030_),
    .C(_1031_),
    .D(_1036_),
    .X(_2064_));
 sky130_fd_sc_hd__and3_2 _5251_ (.A(net185),
    .B(_1159_),
    .C(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__and3b_1 _5252_ (.A_N(net178),
    .B(_1034_),
    .C(net185),
    .X(_2066_));
 sky130_fd_sc_hd__and2_2 _5253_ (.A(_2062_),
    .B(_2066_),
    .X(_2067_));
 sky130_fd_sc_hd__and3_1 _5254_ (.A(net106),
    .B(_2064_),
    .C(_2066_),
    .X(_2068_));
 sky130_fd_sc_hd__a221o_1 _5255_ (.A1(\core_0.execute.sreg_irq_pc.o_d[0] ),
    .A2(_2065_),
    .B1(_2067_),
    .B2(\core_0.execute.sreg_scratch.o_d[0] ),
    .C1(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__and3_2 _5256_ (.A(_1033_),
    .B(_1159_),
    .C(_2061_),
    .X(_2070_));
 sky130_fd_sc_hd__and2_1 _5257_ (.A(net187),
    .B(net186),
    .X(_2071_));
 sky130_fd_sc_hd__and3_1 _5258_ (.A(_1033_),
    .B(_1159_),
    .C(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__a22o_1 _5259_ (.A1(\core_0.execute.sreg_irq_flags.o_d[0] ),
    .A2(_2070_),
    .B1(_2072_),
    .B2(\core_0.execute.pc_high_buff_out[0] ),
    .X(_2073_));
 sky130_fd_sc_hd__and3_1 _5260_ (.A(_1032_),
    .B(_1035_),
    .C(_2071_),
    .X(_2074_));
 sky130_fd_sc_hd__clkbuf_4 _5261_ (.A(_2074_),
    .X(_2075_));
 sky130_fd_sc_hd__and4b_4 _5262_ (.A_N(net186),
    .B(_1032_),
    .C(_1159_),
    .D(net187),
    .X(_2076_));
 sky130_fd_sc_hd__a22o_1 _5263_ (.A1(\core_0.execute.pc_high_out[0] ),
    .A2(_2075_),
    .B1(_2076_),
    .B2(net1),
    .X(_2077_));
 sky130_fd_sc_hd__a22o_1 _5264_ (.A1(net72),
    .A2(_1037_),
    .B1(_1161_),
    .B2(\core_0.execute.sreg_priv_control.o_d[0] ),
    .X(_2078_));
 sky130_fd_sc_hd__and3_2 _5265_ (.A(_1033_),
    .B(_1035_),
    .C(_2061_),
    .X(_2079_));
 sky130_fd_sc_hd__nand2_1 _5266_ (.A(\core_0.execute.alu_flag_reg.o_d[0] ),
    .B(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__or4b_2 _5267_ (.A(_2073_),
    .B(_2077_),
    .C(_2078_),
    .D_N(_2080_),
    .X(_2081_));
 sky130_fd_sc_hd__clkinv_4 _5268_ (.A(\core_0.dec_sreg_jal_over ),
    .Y(_2082_));
 sky130_fd_sc_hd__o32ai_4 _5269_ (.A1(_2063_),
    .A2(_2069_),
    .A3(_2081_),
    .B1(_2082_),
    .B2(net72),
    .Y(_2083_));
 sky130_fd_sc_hd__a21o_1 _5270_ (.A1(_1789_),
    .A2(_2083_),
    .B1(_1792_),
    .X(_2084_));
 sky130_fd_sc_hd__xnor2_1 _5271_ (.A(\core_0.dec_sreg_jal_over ),
    .B(_2084_),
    .Y(_2085_));
 sky130_fd_sc_hd__or2_4 _5272_ (.A(\core_0.dec_sreg_jal_over ),
    .B(\core_0.dec_sreg_load ),
    .X(_2086_));
 sky130_fd_sc_hd__clkbuf_4 _5273_ (.A(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__mux2_1 _5274_ (.A0(_1787_),
    .A1(_2085_),
    .S(_2087_),
    .X(_2088_));
 sky130_fd_sc_hd__buf_4 _5275_ (.A(\core_0.dec_mem_access ),
    .X(_2089_));
 sky130_fd_sc_hd__mux2_1 _5276_ (.A0(_2088_),
    .A1(net194),
    .S(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__mux2_1 _5277_ (.A0(_2090_),
    .A1(\core_0.ew_data[0] ),
    .S(_2044_),
    .X(_2091_));
 sky130_fd_sc_hd__clkbuf_1 _5278_ (.A(_2091_),
    .X(_0229_));
 sky130_fd_sc_hd__a21bo_1 _5279_ (.A1(\core_0.execute.alu_mul_div.div_res[1] ),
    .A2(_1696_),
    .B1_N(_0741_),
    .X(_2092_));
 sky130_fd_sc_hd__mux2_1 _5280_ (.A0(_2010_),
    .A1(_1980_),
    .S(_1422_),
    .X(_2093_));
 sky130_fd_sc_hd__or2_1 _5281_ (.A(_1998_),
    .B(_2093_),
    .X(_2094_));
 sky130_fd_sc_hd__xnor2_1 _5282_ (.A(_1703_),
    .B(_1966_),
    .Y(_2095_));
 sky130_fd_sc_hd__or3b_2 _5283_ (.A(_2095_),
    .B(_1985_),
    .C_N(_1707_),
    .X(_2096_));
 sky130_fd_sc_hd__nor2_2 _5284_ (.A(_1701_),
    .B(_1752_),
    .Y(_2097_));
 sky130_fd_sc_hd__nand2_1 _5285_ (.A(_1751_),
    .B(_2097_),
    .Y(_2098_));
 sky130_fd_sc_hd__nor4_4 _5286_ (.A(_1493_),
    .B(_1344_),
    .C(_1482_),
    .D(_1391_),
    .Y(_2099_));
 sky130_fd_sc_hd__mux2_1 _5287_ (.A0(_1601_),
    .A1(_1841_),
    .S(_1729_),
    .X(_2100_));
 sky130_fd_sc_hd__and3b_1 _5288_ (.A_N(_1733_),
    .B(_2099_),
    .C(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__nor3_4 _5289_ (.A(_1541_),
    .B(_1733_),
    .C(_1734_),
    .Y(_2102_));
 sky130_fd_sc_hd__nor2_2 _5290_ (.A(_1738_),
    .B(_1764_),
    .Y(_2103_));
 sky130_fd_sc_hd__a22oi_2 _5291_ (.A1(_1739_),
    .A2(_2101_),
    .B1(_2102_),
    .B2(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__mux2_1 _5292_ (.A0(_1756_),
    .A1(_1914_),
    .S(_1421_),
    .X(_2105_));
 sky130_fd_sc_hd__mux2_1 _5293_ (.A0(_1550_),
    .A1(_1557_),
    .S(_1729_),
    .X(_2106_));
 sky130_fd_sc_hd__or4b_1 _5294_ (.A(_1724_),
    .B(_1733_),
    .C(_1734_),
    .D_N(_2106_),
    .X(_2107_));
 sky130_fd_sc_hd__o31a_1 _5295_ (.A1(_1739_),
    .A2(_1728_),
    .A3(_2105_),
    .B1(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__mux2_1 _5296_ (.A0(_2104_),
    .A1(_2108_),
    .S(_1431_),
    .X(_2109_));
 sky130_fd_sc_hd__and2b_1 _5297_ (.A_N(_1946_),
    .B(_1943_),
    .X(_2110_));
 sky130_fd_sc_hd__or2_1 _5298_ (.A(_2110_),
    .B(_1944_),
    .X(_2111_));
 sky130_fd_sc_hd__a21oi_1 _5299_ (.A1(_2110_),
    .A2(_1944_),
    .B1(_1773_),
    .Y(_2112_));
 sky130_fd_sc_hd__nor2_1 _5300_ (.A(\core_0.decode.oc_alu_mode[3] ),
    .B(_1775_),
    .Y(_2113_));
 sky130_fd_sc_hd__nor2_1 _5301_ (.A(_1624_),
    .B(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__a221o_1 _5302_ (.A1(\core_0.decode.oc_alu_mode[7] ),
    .A2(_1725_),
    .B1(_1943_),
    .B2(\core_0.decode.oc_alu_mode[9] ),
    .C1(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__a221o_1 _5303_ (.A1(\core_0.decode.oc_alu_mode[2] ),
    .A2(_1946_),
    .B1(_2110_),
    .B2(\core_0.decode.oc_alu_mode[6] ),
    .C1(_2115_),
    .X(_2116_));
 sky130_fd_sc_hd__a21oi_1 _5304_ (.A1(_1885_),
    .A2(_1884_),
    .B1(_1739_),
    .Y(_2117_));
 sky130_fd_sc_hd__a31o_1 _5305_ (.A1(_1739_),
    .A2(_1885_),
    .A3(_1884_),
    .B1(_1774_),
    .X(_2118_));
 sky130_fd_sc_hd__nor2_1 _5306_ (.A(_2117_),
    .B(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__a211oi_1 _5307_ (.A1(_2111_),
    .A2(_2112_),
    .B1(_2116_),
    .C1(_2119_),
    .Y(_2120_));
 sky130_fd_sc_hd__mux2_1 _5308_ (.A0(_1571_),
    .A1(_1579_),
    .S(_1729_),
    .X(_2121_));
 sky130_fd_sc_hd__or4b_1 _5309_ (.A(_1738_),
    .B(_1733_),
    .C(_1734_),
    .D_N(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__mux2_1 _5310_ (.A0(_1654_),
    .A1(_1661_),
    .S(_1421_),
    .X(_2123_));
 sky130_fd_sc_hd__or4b_1 _5311_ (.A(_1724_),
    .B(_1733_),
    .C(_1734_),
    .D_N(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__a21o_1 _5312_ (.A1(_2122_),
    .A2(_2124_),
    .B1(_1431_),
    .X(_2125_));
 sky130_fd_sc_hd__or2_2 _5313_ (.A(_1421_),
    .B(_1677_),
    .X(_2126_));
 sky130_fd_sc_hd__o21ai_1 _5314_ (.A1(_1764_),
    .A2(_1670_),
    .B1(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__nor2_2 _5315_ (.A(_1422_),
    .B(_1633_),
    .Y(_2128_));
 sky130_fd_sc_hd__a211o_1 _5316_ (.A1(_1422_),
    .A2(_1732_),
    .B1(_2128_),
    .C1(_1725_),
    .X(_2129_));
 sky130_fd_sc_hd__o2111ai_1 _5317_ (.A1(_1739_),
    .A2(_2127_),
    .B1(_2129_),
    .C1(_1735_),
    .D1(_1431_),
    .Y(_2130_));
 sky130_fd_sc_hd__nand2_4 _5318_ (.A(_1371_),
    .B(_2097_),
    .Y(_2131_));
 sky130_fd_sc_hd__a21o_1 _5319_ (.A1(_2125_),
    .A2(_2130_),
    .B1(_2131_),
    .X(_2132_));
 sky130_fd_sc_hd__o211a_1 _5320_ (.A1(_2098_),
    .A2(_2109_),
    .B1(_2120_),
    .C1(_2132_),
    .X(_2133_));
 sky130_fd_sc_hd__o21ai_2 _5321_ (.A1(_2094_),
    .A2(_2096_),
    .B1(_2133_),
    .Y(_2134_));
 sky130_fd_sc_hd__clkbuf_4 _5322_ (.A(\core_0.execute.alu_mul_div.i_mul ),
    .X(_2135_));
 sky130_fd_sc_hd__a21o_1 _5323_ (.A1(_2135_),
    .A2(\core_0.execute.alu_mul_div.mul_res[1] ),
    .B1(_0988_),
    .X(_2136_));
 sky130_fd_sc_hd__a21o_1 _5324_ (.A1(_1784_),
    .A2(_2134_),
    .B1(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__a22o_2 _5325_ (.A1(\core_0.execute.alu_mul_div.div_cur[1] ),
    .A2(\core_0.execute.alu_mul_div.i_mod ),
    .B1(_2092_),
    .B2(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__nor2_1 _5326_ (.A(net79),
    .B(_2082_),
    .Y(_2139_));
 sky130_fd_sc_hd__a22o_1 _5327_ (.A1(\core_0.execute.sreg_irq_flags.o_d[1] ),
    .A2(_2070_),
    .B1(_2079_),
    .B2(\core_0.execute.alu_flag_reg.o_d[1] ),
    .X(_2140_));
 sky130_fd_sc_hd__and3_1 _5328_ (.A(\core_0.execute.trap_flag ),
    .B(_2064_),
    .C(_2066_),
    .X(_2141_));
 sky130_fd_sc_hd__and3_1 _5329_ (.A(\core_0.execute.sreg_scratch.o_d[1] ),
    .B(_2062_),
    .C(_2066_),
    .X(_2142_));
 sky130_fd_sc_hd__a2111o_1 _5330_ (.A1(\core_0.execute.sreg_irq_pc.o_d[1] ),
    .A2(_2065_),
    .B1(_2141_),
    .C1(_2142_),
    .D1(\core_0.dec_sreg_jal_over ),
    .X(_2143_));
 sky130_fd_sc_hd__and4_1 _5331_ (.A(\core_0.execute.pc_high_out[1] ),
    .B(_1033_),
    .C(_1035_),
    .D(_2071_),
    .X(_2144_));
 sky130_fd_sc_hd__and4_1 _5332_ (.A(\core_0.execute.pc_high_buff_out[1] ),
    .B(_1033_),
    .C(_1159_),
    .D(_2071_),
    .X(_2145_));
 sky130_fd_sc_hd__and4_1 _5333_ (.A(net79),
    .B(_1033_),
    .C(_1035_),
    .D(_1036_),
    .X(_2146_));
 sky130_fd_sc_hd__a2111o_1 _5334_ (.A1(net8),
    .A2(_2076_),
    .B1(_2144_),
    .C1(_2145_),
    .D1(_2146_),
    .X(_2147_));
 sky130_fd_sc_hd__a2111oi_1 _5335_ (.A1(\core_0.execute.sreg_data_page ),
    .A2(_1161_),
    .B1(_2140_),
    .C1(_2143_),
    .D1(_2147_),
    .Y(_2148_));
 sky130_fd_sc_hd__nand2_1 _5336_ (.A(\core_0.execute.sreg_irq_pc.o_d[1] ),
    .B(\core_0.dec_sreg_irt ),
    .Y(_2149_));
 sky130_fd_sc_hd__o31a_1 _5337_ (.A1(\core_0.dec_sreg_irt ),
    .A2(_2139_),
    .A3(_2148_),
    .B1(_2149_),
    .X(_2150_));
 sky130_fd_sc_hd__a2111oi_4 _5338_ (.A1(_1788_),
    .A2(_2083_),
    .B1(_2150_),
    .C1(_2082_),
    .D1(_1792_),
    .Y(_2151_));
 sky130_fd_sc_hd__clkbuf_4 _5339_ (.A(_2082_),
    .X(_2152_));
 sky130_fd_sc_hd__o21ai_1 _5340_ (.A1(_2152_),
    .A2(_2084_),
    .B1(_2150_),
    .Y(_2153_));
 sky130_fd_sc_hd__and2b_1 _5341_ (.A_N(_2151_),
    .B(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__mux2_1 _5342_ (.A0(_2138_),
    .A1(_2154_),
    .S(_2087_),
    .X(_2155_));
 sky130_fd_sc_hd__mux2_1 _5343_ (.A0(_2155_),
    .A1(net201),
    .S(_2089_),
    .X(_2156_));
 sky130_fd_sc_hd__mux2_1 _5344_ (.A0(_2156_),
    .A1(\core_0.ew_data[1] ),
    .S(_2044_),
    .X(_2157_));
 sky130_fd_sc_hd__clkbuf_1 _5345_ (.A(_2157_),
    .X(_0230_));
 sky130_fd_sc_hd__nor2_1 _5346_ (.A(\core_0.dec_sreg_jal_over ),
    .B(\core_0.dec_sreg_load ),
    .Y(_2158_));
 sky130_fd_sc_hd__clkbuf_4 _5347_ (.A(_2158_),
    .X(_2159_));
 sky130_fd_sc_hd__a21bo_1 _5348_ (.A1(\core_0.execute.alu_mul_div.div_res[2] ),
    .A2(_1697_),
    .B1_N(_1411_),
    .X(_2160_));
 sky130_fd_sc_hd__mux2_1 _5349_ (.A0(_1979_),
    .A1(_1980_),
    .S(_1764_),
    .X(_2161_));
 sky130_fd_sc_hd__o2bb2a_1 _5350_ (.A1_N(_1723_),
    .A2_N(_2103_),
    .B1(_2161_),
    .B2(_1998_),
    .X(_2162_));
 sky130_fd_sc_hd__a21oi_1 _5351_ (.A1(_1943_),
    .A2(_1944_),
    .B1(_1946_),
    .Y(_2163_));
 sky130_fd_sc_hd__a221o_1 _5352_ (.A1(\core_0.decode.oc_alu_mode[11] ),
    .A2(_1886_),
    .B1(_2163_),
    .B2(\core_0.decode.oc_alu_mode[4] ),
    .C1(\core_0.decode.oc_alu_mode[6] ),
    .X(_2164_));
 sky130_fd_sc_hd__o22ai_1 _5353_ (.A1(_1774_),
    .A2(_1886_),
    .B1(_2163_),
    .B2(_1773_),
    .Y(_2165_));
 sky130_fd_sc_hd__inv_2 _5354_ (.A(_1945_),
    .Y(_2166_));
 sky130_fd_sc_hd__nand2_1 _5355_ (.A(_1942_),
    .B(_2166_),
    .Y(_2167_));
 sky130_fd_sc_hd__mux2_1 _5356_ (.A0(_2164_),
    .A1(_2165_),
    .S(_2167_),
    .X(_2168_));
 sky130_fd_sc_hd__a2bb2o_1 _5357_ (.A1_N(_1633_),
    .A2_N(_2113_),
    .B1(\core_0.decode.oc_alu_mode[7] ),
    .B2(_1741_),
    .X(_2169_));
 sky130_fd_sc_hd__a221o_1 _5358_ (.A1(\core_0.decode.oc_alu_mode[9] ),
    .A2(_1942_),
    .B1(_1945_),
    .B2(\core_0.decode.oc_alu_mode[2] ),
    .C1(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__nor2_1 _5359_ (.A(_2168_),
    .B(_2170_),
    .Y(_2171_));
 sky130_fd_sc_hd__mux2_1 _5360_ (.A0(_1920_),
    .A1(_1914_),
    .S(_1729_),
    .X(_2172_));
 sky130_fd_sc_hd__mux2_1 _5361_ (.A0(_1758_),
    .A1(_2172_),
    .S(_1739_),
    .X(_2173_));
 sky130_fd_sc_hd__or4_1 _5362_ (.A(_1374_),
    .B(_1725_),
    .C(_1727_),
    .D(_1755_),
    .X(_2174_));
 sky130_fd_sc_hd__o31a_1 _5363_ (.A1(_1741_),
    .A2(_1728_),
    .A3(_2173_),
    .B1(_2174_),
    .X(_2175_));
 sky130_fd_sc_hd__mux2_1 _5364_ (.A0(_1549_),
    .A1(_1579_),
    .S(_1421_),
    .X(_2176_));
 sky130_fd_sc_hd__or4b_1 _5365_ (.A(_1738_),
    .B(_1726_),
    .C(_1734_),
    .D_N(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__o31a_1 _5366_ (.A1(_1725_),
    .A2(_1727_),
    .A3(_1747_),
    .B1(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__o31a_1 _5367_ (.A1(_1733_),
    .A2(_1734_),
    .A3(_1730_),
    .B1(_1738_),
    .X(_2179_));
 sky130_fd_sc_hd__o31a_1 _5368_ (.A1(_1733_),
    .A2(_1734_),
    .A3(_1744_),
    .B1(_1724_),
    .X(_2180_));
 sky130_fd_sc_hd__or3_1 _5369_ (.A(_1698_),
    .B(_2179_),
    .C(_2180_),
    .X(_2181_));
 sky130_fd_sc_hd__o211a_1 _5370_ (.A1(_1431_),
    .A2(_2178_),
    .B1(_2181_),
    .C1(_1371_),
    .X(_2182_));
 sky130_fd_sc_hd__a211o_1 _5371_ (.A1(_1751_),
    .A2(_2175_),
    .B1(_2182_),
    .C1(_1753_),
    .X(_2183_));
 sky130_fd_sc_hd__o211a_1 _5372_ (.A1(_2096_),
    .A2(_2162_),
    .B1(_2171_),
    .C1(_2183_),
    .X(_2184_));
 sky130_fd_sc_hd__nor2_1 _5373_ (.A(_2135_),
    .B(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__a211o_1 _5374_ (.A1(_0955_),
    .A2(\core_0.execute.alu_mul_div.mul_res[2] ),
    .B1(_2185_),
    .C1(_0989_),
    .X(_2186_));
 sky130_fd_sc_hd__a22o_2 _5375_ (.A1(\core_0.execute.alu_mul_div.div_cur[2] ),
    .A2(_0960_),
    .B1(_2160_),
    .B2(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__or2_1 _5376_ (.A(\core_0.dec_sreg_jal_over ),
    .B(_1037_),
    .X(_2188_));
 sky130_fd_sc_hd__and2_1 _5377_ (.A(net80),
    .B(_2188_),
    .X(_2189_));
 sky130_fd_sc_hd__a22o_1 _5378_ (.A1(\core_0.execute.pc_high_out[2] ),
    .A2(_2075_),
    .B1(_2079_),
    .B2(\core_0.execute.alu_flag_reg.o_d[2] ),
    .X(_2190_));
 sky130_fd_sc_hd__a221o_1 _5379_ (.A1(\core_0.execute.irq_en ),
    .A2(_1161_),
    .B1(_2070_),
    .B2(\core_0.execute.sreg_irq_flags.o_d[2] ),
    .C1(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__and4_1 _5380_ (.A(net187),
    .B(net186),
    .C(_1033_),
    .D(_1159_),
    .X(_2192_));
 sky130_fd_sc_hd__and4b_4 _5381_ (.A_N(net186),
    .B(_1033_),
    .C(_1159_),
    .D(net187),
    .X(_2193_));
 sky130_fd_sc_hd__and3_1 _5382_ (.A(net105),
    .B(_2064_),
    .C(_2066_),
    .X(_2194_));
 sky130_fd_sc_hd__a221o_1 _5383_ (.A1(\core_0.execute.sreg_irq_pc.o_d[2] ),
    .A2(_2065_),
    .B1(_2067_),
    .B2(\core_0.execute.sreg_scratch.o_d[2] ),
    .C1(_2194_),
    .X(_2195_));
 sky130_fd_sc_hd__a221o_1 _5384_ (.A1(\core_0.execute.pc_high_buff_out[2] ),
    .A2(_2192_),
    .B1(_2193_),
    .B2(net9),
    .C1(_2195_),
    .X(_2196_));
 sky130_fd_sc_hd__o21a_1 _5385_ (.A1(_2191_),
    .A2(_2196_),
    .B1(_2082_),
    .X(_2197_));
 sky130_fd_sc_hd__or2_1 _5386_ (.A(\core_0.execute.sreg_irq_pc.o_d[2] ),
    .B(_1788_),
    .X(_2198_));
 sky130_fd_sc_hd__o31a_2 _5387_ (.A1(\core_0.dec_sreg_irt ),
    .A2(_2189_),
    .A3(_2197_),
    .B1(_2198_),
    .X(_2199_));
 sky130_fd_sc_hd__nand2_1 _5388_ (.A(_2151_),
    .B(_2199_),
    .Y(_2200_));
 sky130_fd_sc_hd__o21a_1 _5389_ (.A1(_2151_),
    .A2(_2199_),
    .B1(_2086_),
    .X(_2201_));
 sky130_fd_sc_hd__a22o_1 _5390_ (.A1(_2159_),
    .A2(_2187_),
    .B1(_2200_),
    .B2(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__mux2_1 _5391_ (.A0(_2202_),
    .A1(net202),
    .S(_2089_),
    .X(_2203_));
 sky130_fd_sc_hd__mux2_1 _5392_ (.A0(_2203_),
    .A1(\core_0.ew_data[2] ),
    .S(_2044_),
    .X(_2204_));
 sky130_fd_sc_hd__clkbuf_1 _5393_ (.A(_2204_),
    .X(_0231_));
 sky130_fd_sc_hd__and2_2 _5394_ (.A(\core_0.execute.sreg_irq_pc.o_d[3] ),
    .B(\core_0.dec_sreg_irt ),
    .X(_2205_));
 sky130_fd_sc_hd__a22o_1 _5395_ (.A1(net81),
    .A2(_1037_),
    .B1(_2070_),
    .B2(\core_0.execute.sreg_irq_flags.o_d[3] ),
    .X(_2206_));
 sky130_fd_sc_hd__a221o_1 _5396_ (.A1(\core_0.execute.sreg_irq_pc.o_d[3] ),
    .A2(_2065_),
    .B1(_2067_),
    .B2(\core_0.execute.sreg_scratch.o_d[3] ),
    .C1(\core_0.dec_sreg_jal_over ),
    .X(_2207_));
 sky130_fd_sc_hd__a22o_1 _5397_ (.A1(\core_0.execute.pc_high_out[3] ),
    .A2(_2075_),
    .B1(_2079_),
    .B2(\core_0.execute.alu_flag_reg.o_d[3] ),
    .X(_2208_));
 sky130_fd_sc_hd__a221o_1 _5398_ (.A1(\core_0.execute.pc_high_buff_out[3] ),
    .A2(_2072_),
    .B1(_2076_),
    .B2(net10),
    .C1(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__a211o_1 _5399_ (.A1(\core_0.execute.sreg_long_ptr_en ),
    .A2(_1161_),
    .B1(_2207_),
    .C1(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__o221a_2 _5400_ (.A1(net81),
    .A2(_2082_),
    .B1(_2206_),
    .B2(_2210_),
    .C1(_1788_),
    .X(_2211_));
 sky130_fd_sc_hd__a211oi_1 _5401_ (.A1(_2151_),
    .A2(_2199_),
    .B1(_2205_),
    .C1(_2211_),
    .Y(_2212_));
 sky130_fd_sc_hd__o211ai_4 _5402_ (.A1(_2205_),
    .A2(_2211_),
    .B1(_2151_),
    .C1(_2199_),
    .Y(_2213_));
 sky130_fd_sc_hd__nand2_1 _5403_ (.A(_2086_),
    .B(_2213_),
    .Y(_2214_));
 sky130_fd_sc_hd__a21bo_1 _5404_ (.A1(\core_0.execute.alu_mul_div.div_res[3] ),
    .A2(_1697_),
    .B1_N(_1411_),
    .X(_2215_));
 sky130_fd_sc_hd__or4_1 _5405_ (.A(_1724_),
    .B(_1733_),
    .C(_1734_),
    .D(_2105_),
    .X(_2216_));
 sky130_fd_sc_hd__a21bo_2 _5406_ (.A1(_1725_),
    .A2(_2101_),
    .B1_N(_2216_),
    .X(_2217_));
 sky130_fd_sc_hd__and3_1 _5407_ (.A(_1741_),
    .B(_1983_),
    .C(_2102_),
    .X(_2218_));
 sky130_fd_sc_hd__a211o_1 _5408_ (.A1(_1431_),
    .A2(_2217_),
    .B1(_2218_),
    .C1(_1371_),
    .X(_2219_));
 sky130_fd_sc_hd__and4b_1 _5409_ (.A_N(_1733_),
    .B(_2106_),
    .C(_2099_),
    .D(_1725_),
    .X(_2220_));
 sky130_fd_sc_hd__a31o_1 _5410_ (.A1(_1739_),
    .A2(_1735_),
    .A3(_2121_),
    .B1(_2220_),
    .X(_2221_));
 sky130_fd_sc_hd__mux2_1 _5411_ (.A0(_2123_),
    .A1(_2127_),
    .S(_1739_),
    .X(_2222_));
 sky130_fd_sc_hd__nor2_1 _5412_ (.A(_1741_),
    .B(_1728_),
    .Y(_2223_));
 sky130_fd_sc_hd__a221o_1 _5413_ (.A1(_1749_),
    .A2(_2221_),
    .B1(_2222_),
    .B2(_2223_),
    .C1(_1751_),
    .X(_2224_));
 sky130_fd_sc_hd__nand3_2 _5414_ (.A(_2097_),
    .B(_2219_),
    .C(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__a21oi_1 _5415_ (.A1(_1881_),
    .A2(_1886_),
    .B1(_1887_),
    .Y(_2226_));
 sky130_fd_sc_hd__xnor2_1 _5416_ (.A(_1890_),
    .B(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__mux4_1 _5417_ (.A0(_2010_),
    .A1(_1979_),
    .A2(_1980_),
    .A3(_1978_),
    .S0(_1975_),
    .S1(_1422_),
    .X(_2228_));
 sky130_fd_sc_hd__inv_2 _5418_ (.A(\core_0.decode.oc_alu_mode[6] ),
    .Y(_2229_));
 sky130_fd_sc_hd__nor2_1 _5419_ (.A(_2229_),
    .B(_1888_),
    .Y(_2230_));
 sky130_fd_sc_hd__a221o_4 _5420_ (.A1(net97),
    .A2(_1563_),
    .B1(_1665_),
    .B2(_0715_),
    .C1(_1669_),
    .X(_2231_));
 sky130_fd_sc_hd__a221o_1 _5421_ (.A1(\core_0.decode.oc_alu_mode[7] ),
    .A2(_1703_),
    .B1(_2231_),
    .B2(_1776_),
    .C1(\core_0.decode.oc_alu_mode[9] ),
    .X(_2232_));
 sky130_fd_sc_hd__a211o_1 _5422_ (.A1(\core_0.decode.oc_alu_mode[2] ),
    .A2(_1888_),
    .B1(_2230_),
    .C1(_2232_),
    .X(_2233_));
 sky130_fd_sc_hd__a31o_1 _5423_ (.A1(_1890_),
    .A2(_1942_),
    .A3(_1947_),
    .B1(_1773_),
    .X(_2234_));
 sky130_fd_sc_hd__a21oi_1 _5424_ (.A1(_1942_),
    .A2(_1947_),
    .B1(_1890_),
    .Y(_2235_));
 sky130_fd_sc_hd__o2bb2a_1 _5425_ (.A1_N(_1889_),
    .A2_N(_2233_),
    .B1(_2234_),
    .B2(_2235_),
    .X(_2236_));
 sky130_fd_sc_hd__o221a_1 _5426_ (.A1(_1774_),
    .A2(_2227_),
    .B1(_2228_),
    .B2(_2096_),
    .C1(_2236_),
    .X(_2237_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(_2225_),
    .B(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__a21o_1 _5428_ (.A1(_2135_),
    .A2(\core_0.execute.alu_mul_div.mul_res[3] ),
    .B1(_0988_),
    .X(_2239_));
 sky130_fd_sc_hd__a21o_1 _5429_ (.A1(_1784_),
    .A2(_2238_),
    .B1(_2239_),
    .X(_2240_));
 sky130_fd_sc_hd__a22o_2 _5430_ (.A1(\core_0.execute.alu_mul_div.div_cur[3] ),
    .A2(_0960_),
    .B1(_2215_),
    .B2(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__a2bb2o_1 _5431_ (.A1_N(_2212_),
    .A2_N(_2214_),
    .B1(_2159_),
    .B2(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__mux2_1 _5432_ (.A0(_2242_),
    .A1(net203),
    .S(_2089_),
    .X(_2243_));
 sky130_fd_sc_hd__mux2_1 _5433_ (.A0(_2243_),
    .A1(\core_0.ew_data[3] ),
    .S(_2044_),
    .X(_2244_));
 sky130_fd_sc_hd__clkbuf_1 _5434_ (.A(_2244_),
    .X(_0232_));
 sky130_fd_sc_hd__a21bo_1 _5435_ (.A1(\core_0.execute.alu_mul_div.div_res[4] ),
    .A2(_1697_),
    .B1_N(_1411_),
    .X(_2245_));
 sky130_fd_sc_hd__nand2_2 _5436_ (.A(_1707_),
    .B(_1967_),
    .Y(_2246_));
 sky130_fd_sc_hd__nor2_1 _5437_ (.A(_1431_),
    .B(_1699_),
    .Y(_2247_));
 sky130_fd_sc_hd__o2bb2a_1 _5438_ (.A1_N(_1723_),
    .A2_N(_2247_),
    .B1(_1982_),
    .B2(_1985_),
    .X(_2248_));
 sky130_fd_sc_hd__nor2_1 _5439_ (.A(_2246_),
    .B(_2248_),
    .Y(_2249_));
 sky130_fd_sc_hd__mux2_1 _5440_ (.A0(_1895_),
    .A1(_1897_),
    .S(_1891_),
    .X(_2250_));
 sky130_fd_sc_hd__nor2_1 _5441_ (.A(_1774_),
    .B(_2250_),
    .Y(_2251_));
 sky130_fd_sc_hd__nand2_1 _5442_ (.A(_1895_),
    .B(_1948_),
    .Y(_2252_));
 sky130_fd_sc_hd__or2_1 _5443_ (.A(_1895_),
    .B(_1948_),
    .X(_2253_));
 sky130_fd_sc_hd__and3_1 _5444_ (.A(\core_0.decode.oc_alu_mode[4] ),
    .B(_2252_),
    .C(_2253_),
    .X(_2254_));
 sky130_fd_sc_hd__o31ai_1 _5445_ (.A1(_1741_),
    .A2(_1728_),
    .A3(_1748_),
    .B1(_1371_),
    .Y(_2255_));
 sky130_fd_sc_hd__a31o_1 _5446_ (.A1(_1749_),
    .A2(_1735_),
    .A3(_1760_),
    .B1(_2255_),
    .X(_2256_));
 sky130_fd_sc_hd__or3_1 _5447_ (.A(_1741_),
    .B(_1728_),
    .C(_1759_),
    .X(_2257_));
 sky130_fd_sc_hd__nand2_1 _5448_ (.A(_1751_),
    .B(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__nor2_1 _5449_ (.A(_1677_),
    .B(_2113_),
    .Y(_2259_));
 sky130_fd_sc_hd__a221o_1 _5450_ (.A1(\core_0.decode.oc_alu_mode[7] ),
    .A2(_1701_),
    .B1(_1893_),
    .B2(\core_0.decode.oc_alu_mode[9] ),
    .C1(_2259_),
    .X(_2260_));
 sky130_fd_sc_hd__a221o_1 _5451_ (.A1(\core_0.decode.oc_alu_mode[2] ),
    .A2(_1892_),
    .B1(_1895_),
    .B2(\core_0.decode.oc_alu_mode[6] ),
    .C1(_2260_),
    .X(_2261_));
 sky130_fd_sc_hd__a31o_1 _5452_ (.A1(_2097_),
    .A2(_2256_),
    .A3(_2258_),
    .B1(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__or4_2 _5453_ (.A(_2249_),
    .B(_2251_),
    .C(_2254_),
    .D(_2262_),
    .X(_2263_));
 sky130_fd_sc_hd__a21o_1 _5454_ (.A1(_2135_),
    .A2(\core_0.execute.alu_mul_div.mul_res[4] ),
    .B1(_0988_),
    .X(_2264_));
 sky130_fd_sc_hd__a21o_1 _5455_ (.A1(_1784_),
    .A2(_2263_),
    .B1(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__a22o_2 _5456_ (.A1(\core_0.execute.alu_mul_div.div_cur[4] ),
    .A2(_0960_),
    .B1(_2245_),
    .B2(_2265_),
    .X(_2266_));
 sky130_fd_sc_hd__a22o_1 _5457_ (.A1(net82),
    .A2(_1037_),
    .B1(_2075_),
    .B2(\core_0.execute.pc_high_out[4] ),
    .X(_2267_));
 sky130_fd_sc_hd__a221o_1 _5458_ (.A1(\core_0.execute.sreg_irq_pc.o_d[4] ),
    .A2(_2065_),
    .B1(_2067_),
    .B2(\core_0.execute.sreg_scratch.o_d[4] ),
    .C1(_2063_),
    .X(_2268_));
 sky130_fd_sc_hd__a221o_1 _5459_ (.A1(\core_0.execute.sreg_priv_control.o_d[4] ),
    .A2(_1161_),
    .B1(_2079_),
    .B2(\core_0.execute.alu_flag_reg.o_d[4] ),
    .C1(_2268_),
    .X(_2269_));
 sky130_fd_sc_hd__a221o_1 _5460_ (.A1(\core_0.execute.pc_high_buff_out[4] ),
    .A2(_2192_),
    .B1(_2193_),
    .B2(net11),
    .C1(_2269_),
    .X(_2270_));
 sky130_fd_sc_hd__a211oi_1 _5461_ (.A1(\core_0.execute.sreg_irq_flags.o_d[4] ),
    .A2(_2070_),
    .B1(_2267_),
    .C1(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__nor2_1 _5462_ (.A(net82),
    .B(_2082_),
    .Y(_2272_));
 sky130_fd_sc_hd__nand2_1 _5463_ (.A(\core_0.execute.sreg_irq_pc.o_d[4] ),
    .B(\core_0.dec_sreg_irt ),
    .Y(_2273_));
 sky130_fd_sc_hd__o31a_2 _5464_ (.A1(\core_0.dec_sreg_irt ),
    .A2(_2271_),
    .A3(_2272_),
    .B1(_2273_),
    .X(_2274_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(_2213_),
    .B(_2274_),
    .Y(_2275_));
 sky130_fd_sc_hd__o21a_1 _5466_ (.A1(_2213_),
    .A2(_2274_),
    .B1(_2086_),
    .X(_2276_));
 sky130_fd_sc_hd__a22o_1 _5467_ (.A1(_2159_),
    .A2(_2266_),
    .B1(_2275_),
    .B2(_2276_),
    .X(_2277_));
 sky130_fd_sc_hd__mux2_1 _5468_ (.A0(_2277_),
    .A1(net204),
    .S(_2089_),
    .X(_2278_));
 sky130_fd_sc_hd__mux2_1 _5469_ (.A0(_2278_),
    .A1(\core_0.ew_data[4] ),
    .S(_2044_),
    .X(_2279_));
 sky130_fd_sc_hd__clkbuf_1 _5470_ (.A(_2279_),
    .X(_0233_));
 sky130_fd_sc_hd__a21bo_1 _5471_ (.A1(\core_0.execute.alu_mul_div.div_res[5] ),
    .A2(_1696_),
    .B1_N(_0741_),
    .X(_2280_));
 sky130_fd_sc_hd__mux4_1 _5472_ (.A0(_1969_),
    .A1(_1977_),
    .A2(_1978_),
    .A3(_1979_),
    .S0(_2002_),
    .S1(_1998_),
    .X(_2281_));
 sky130_fd_sc_hd__mux2_1 _5473_ (.A0(_2094_),
    .A1(_2281_),
    .S(_1988_),
    .X(_2282_));
 sky130_fd_sc_hd__a21oi_1 _5474_ (.A1(_1891_),
    .A2(_1896_),
    .B1(_1895_),
    .Y(_2283_));
 sky130_fd_sc_hd__xnor2_1 _5475_ (.A(_1880_),
    .B(_2283_),
    .Y(_2284_));
 sky130_fd_sc_hd__a21o_1 _5476_ (.A1(_1895_),
    .A2(_1948_),
    .B1(_1892_),
    .X(_2285_));
 sky130_fd_sc_hd__xnor2_1 _5477_ (.A(_1877_),
    .B(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__a31o_1 _5478_ (.A1(_1374_),
    .A2(_2122_),
    .A3(_2124_),
    .B1(_2131_),
    .X(_2287_));
 sky130_fd_sc_hd__a21oi_1 _5479_ (.A1(_1749_),
    .A2(_2108_),
    .B1(_2287_),
    .Y(_2288_));
 sky130_fd_sc_hd__a221o_1 _5480_ (.A1(\core_0.decode.oc_alu_mode[7] ),
    .A2(_1709_),
    .B1(_1661_),
    .B2(_1776_),
    .C1(\core_0.decode.oc_alu_mode[9] ),
    .X(_2289_));
 sky130_fd_sc_hd__nor2_1 _5481_ (.A(_2229_),
    .B(_1877_),
    .Y(_2290_));
 sky130_fd_sc_hd__a221o_1 _5482_ (.A1(\core_0.decode.oc_alu_mode[2] ),
    .A2(_1952_),
    .B1(_2289_),
    .B2(_1953_),
    .C1(_2290_),
    .X(_2291_));
 sky130_fd_sc_hd__or3_1 _5483_ (.A(_1741_),
    .B(_2098_),
    .C(_2104_),
    .X(_2292_));
 sky130_fd_sc_hd__or3b_1 _5484_ (.A(_2288_),
    .B(_2291_),
    .C_N(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__a221o_1 _5485_ (.A1(\core_0.decode.oc_alu_mode[11] ),
    .A2(_2284_),
    .B1(_2286_),
    .B2(_0962_),
    .C1(_2293_),
    .X(_2294_));
 sky130_fd_sc_hd__o21bai_2 _5486_ (.A1(_2246_),
    .A2(_2282_),
    .B1_N(_2294_),
    .Y(_2295_));
 sky130_fd_sc_hd__a21o_1 _5487_ (.A1(_2135_),
    .A2(\core_0.execute.alu_mul_div.mul_res[5] ),
    .B1(_0988_),
    .X(_2296_));
 sky130_fd_sc_hd__a21o_1 _5488_ (.A1(_1784_),
    .A2(_2295_),
    .B1(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__a22o_4 _5489_ (.A1(\core_0.execute.alu_mul_div.div_cur[5] ),
    .A2(\core_0.execute.alu_mul_div.i_mod ),
    .B1(_2280_),
    .B2(_2297_),
    .X(_2298_));
 sky130_fd_sc_hd__a22o_1 _5490_ (.A1(\core_0.execute.sreg_irq_pc.o_d[5] ),
    .A2(_2065_),
    .B1(_2067_),
    .B2(\core_0.execute.sreg_scratch.o_d[5] ),
    .X(_2299_));
 sky130_fd_sc_hd__a221o_1 _5491_ (.A1(\core_0.execute.sreg_priv_control.o_d[5] ),
    .A2(_1161_),
    .B1(_2075_),
    .B2(\core_0.execute.pc_high_out[5] ),
    .C1(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__a221o_1 _5492_ (.A1(\core_0.execute.pc_high_buff_out[5] ),
    .A2(_2192_),
    .B1(_2193_),
    .B2(net12),
    .C1(_2300_),
    .X(_2301_));
 sky130_fd_sc_hd__a22o_1 _5493_ (.A1(net83),
    .A2(_2188_),
    .B1(_2301_),
    .B2(_2082_),
    .X(_2302_));
 sky130_fd_sc_hd__mux2_1 _5494_ (.A0(\core_0.execute.sreg_irq_pc.o_d[5] ),
    .A1(_2302_),
    .S(_1788_),
    .X(_2303_));
 sky130_fd_sc_hd__nor3b_1 _5495_ (.A(_2213_),
    .B(_2274_),
    .C_N(_2303_),
    .Y(_2304_));
 sky130_fd_sc_hd__o21ba_1 _5496_ (.A1(_2213_),
    .A2(_2274_),
    .B1_N(_2303_),
    .X(_2305_));
 sky130_fd_sc_hd__nor2_1 _5497_ (.A(_2304_),
    .B(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__mux2_1 _5498_ (.A0(_2298_),
    .A1(_2306_),
    .S(_2087_),
    .X(_2307_));
 sky130_fd_sc_hd__mux2_1 _5499_ (.A0(_2307_),
    .A1(net205),
    .S(_2089_),
    .X(_2308_));
 sky130_fd_sc_hd__mux2_1 _5500_ (.A0(_2308_),
    .A1(\core_0.ew_data[5] ),
    .S(_2044_),
    .X(_2309_));
 sky130_fd_sc_hd__clkbuf_1 _5501_ (.A(_2309_),
    .X(_0234_));
 sky130_fd_sc_hd__clkbuf_4 _5502_ (.A(_2188_),
    .X(_2310_));
 sky130_fd_sc_hd__a22o_1 _5503_ (.A1(\core_0.execute.sreg_irq_pc.o_d[6] ),
    .A2(_2065_),
    .B1(_2067_),
    .B2(\core_0.execute.sreg_scratch.o_d[6] ),
    .X(_2311_));
 sky130_fd_sc_hd__a221o_1 _5504_ (.A1(\core_0.execute.sreg_priv_control.o_d[6] ),
    .A2(_1161_),
    .B1(_2075_),
    .B2(\core_0.execute.pc_high_out[6] ),
    .C1(_2311_),
    .X(_2312_));
 sky130_fd_sc_hd__a221o_1 _5505_ (.A1(\core_0.execute.pc_high_buff_out[6] ),
    .A2(_2192_),
    .B1(_2193_),
    .B2(net13),
    .C1(_2312_),
    .X(_2313_));
 sky130_fd_sc_hd__a22o_1 _5506_ (.A1(net84),
    .A2(_2310_),
    .B1(_2313_),
    .B2(_2082_),
    .X(_2314_));
 sky130_fd_sc_hd__mux2_2 _5507_ (.A0(\core_0.execute.sreg_irq_pc.o_d[6] ),
    .A1(_2314_),
    .S(_1788_),
    .X(_2315_));
 sky130_fd_sc_hd__or2_1 _5508_ (.A(_2304_),
    .B(_2315_),
    .X(_2316_));
 sky130_fd_sc_hd__nand2_1 _5509_ (.A(_2304_),
    .B(_2315_),
    .Y(_2317_));
 sky130_fd_sc_hd__a21bo_1 _5510_ (.A1(\core_0.execute.alu_mul_div.div_res[6] ),
    .A2(_1696_),
    .B1_N(_0741_),
    .X(_2318_));
 sky130_fd_sc_hd__o21ba_1 _5511_ (.A1(_1877_),
    .A2(_2252_),
    .B1_N(_1954_),
    .X(_2319_));
 sky130_fd_sc_hd__xnor2_1 _5512_ (.A(_1873_),
    .B(_2319_),
    .Y(_2320_));
 sky130_fd_sc_hd__and2_1 _5513_ (.A(_1707_),
    .B(_1967_),
    .X(_2321_));
 sky130_fd_sc_hd__mux2_1 _5514_ (.A0(_1979_),
    .A1(_1980_),
    .S(_2002_),
    .X(_2322_));
 sky130_fd_sc_hd__a2bb2o_1 _5515_ (.A1_N(_1998_),
    .A2_N(_2322_),
    .B1(_2103_),
    .B2(_1723_),
    .X(_2323_));
 sky130_fd_sc_hd__mux4_2 _5516_ (.A0(_1968_),
    .A1(_1969_),
    .A2(_1977_),
    .A3(_1978_),
    .S0(_1764_),
    .S1(_1981_),
    .X(_2324_));
 sky130_fd_sc_hd__clkinv_2 _5517_ (.A(_2324_),
    .Y(_2325_));
 sky130_fd_sc_hd__mux2_1 _5518_ (.A0(_2323_),
    .A1(_2325_),
    .S(_1988_),
    .X(_2326_));
 sky130_fd_sc_hd__a22o_1 _5519_ (.A1(_0934_),
    .A2(_1357_),
    .B1(_1654_),
    .B2(_1776_),
    .X(_2327_));
 sky130_fd_sc_hd__a221o_1 _5520_ (.A1(_0956_),
    .A2(_1955_),
    .B1(_1873_),
    .B2(_0928_),
    .C1(_2327_),
    .X(_2328_));
 sky130_fd_sc_hd__or4_1 _5521_ (.A(_1749_),
    .B(_1725_),
    .C(_1728_),
    .D(_1755_),
    .X(_2329_));
 sky130_fd_sc_hd__or3_1 _5522_ (.A(_1431_),
    .B(_1728_),
    .C(_2173_),
    .X(_2330_));
 sky130_fd_sc_hd__o211a_1 _5523_ (.A1(_1749_),
    .A2(_2178_),
    .B1(_2330_),
    .C1(_1371_),
    .X(_2331_));
 sky130_fd_sc_hd__a211oi_2 _5524_ (.A1(_1751_),
    .A2(_2329_),
    .B1(_2331_),
    .C1(_1753_),
    .Y(_2332_));
 sky130_fd_sc_hd__a211o_1 _5525_ (.A1(_0998_),
    .A2(_1871_),
    .B1(_2328_),
    .C1(_2332_),
    .X(_2333_));
 sky130_fd_sc_hd__and2_1 _5526_ (.A(_1876_),
    .B(_1899_),
    .X(_2334_));
 sky130_fd_sc_hd__nor2_1 _5527_ (.A(_1774_),
    .B(_2334_),
    .Y(_2335_));
 sky130_fd_sc_hd__o21a_1 _5528_ (.A1(_1876_),
    .A2(_1899_),
    .B1(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__a211o_1 _5529_ (.A1(_2321_),
    .A2(_2326_),
    .B1(_2333_),
    .C1(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__a21oi_2 _5530_ (.A1(_0962_),
    .A2(_2320_),
    .B1(_2337_),
    .Y(_2338_));
 sky130_fd_sc_hd__nor2_1 _5531_ (.A(\core_0.execute.alu_mul_div.i_mul ),
    .B(_2338_),
    .Y(_2339_));
 sky130_fd_sc_hd__a211o_1 _5532_ (.A1(\core_0.execute.alu_mul_div.i_mul ),
    .A2(\core_0.execute.alu_mul_div.mul_res[6] ),
    .B1(_2339_),
    .C1(_0988_),
    .X(_2340_));
 sky130_fd_sc_hd__a22o_4 _5533_ (.A1(\core_0.execute.alu_mul_div.div_cur[6] ),
    .A2(\core_0.execute.alu_mul_div.i_mod ),
    .B1(_2318_),
    .B2(_2340_),
    .X(_2341_));
 sky130_fd_sc_hd__and2_1 _5534_ (.A(_2158_),
    .B(_2341_),
    .X(_2342_));
 sky130_fd_sc_hd__a31o_1 _5535_ (.A1(_2087_),
    .A2(_2316_),
    .A3(_2317_),
    .B1(_2342_),
    .X(_2343_));
 sky130_fd_sc_hd__mux2_1 _5536_ (.A0(_2343_),
    .A1(net206),
    .S(_2089_),
    .X(_2344_));
 sky130_fd_sc_hd__clkbuf_8 _5537_ (.A(_1835_),
    .X(_2345_));
 sky130_fd_sc_hd__mux2_1 _5538_ (.A0(_2344_),
    .A1(\core_0.ew_data[6] ),
    .S(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__clkbuf_1 _5539_ (.A(_2346_),
    .X(_0235_));
 sky130_fd_sc_hd__a21bo_1 _5540_ (.A1(\core_0.execute.alu_mul_div.div_res[7] ),
    .A2(_1697_),
    .B1_N(_1411_),
    .X(_2347_));
 sky130_fd_sc_hd__o21ai_1 _5541_ (.A1(_1875_),
    .A2(_2334_),
    .B1(_1870_),
    .Y(_2348_));
 sky130_fd_sc_hd__or3_1 _5542_ (.A(_1870_),
    .B(_1875_),
    .C(_2334_),
    .X(_2349_));
 sky130_fd_sc_hd__o21ba_1 _5543_ (.A1(_1872_),
    .A2(_2319_),
    .B1_N(_1871_),
    .X(_2350_));
 sky130_fd_sc_hd__xnor2_1 _5544_ (.A(_1867_),
    .B(_2350_),
    .Y(_2351_));
 sky130_fd_sc_hd__mux4_1 _5545_ (.A0(_2010_),
    .A1(_1979_),
    .A2(_1980_),
    .A3(_1978_),
    .S0(_1975_),
    .S1(_1423_),
    .X(_2352_));
 sky130_fd_sc_hd__mux4_1 _5546_ (.A0(_1968_),
    .A1(_1971_),
    .A2(_1977_),
    .A3(_1969_),
    .S0(_1422_),
    .S1(_1998_),
    .X(_2353_));
 sky130_fd_sc_hd__mux2_1 _5547_ (.A0(_2352_),
    .A1(_2353_),
    .S(_1988_),
    .X(_2354_));
 sky130_fd_sc_hd__nor2_1 _5548_ (.A(_1431_),
    .B(_2217_),
    .Y(_2355_));
 sky130_fd_sc_hd__o21ai_2 _5549_ (.A1(_1749_),
    .A2(_2221_),
    .B1(_1754_),
    .Y(_2356_));
 sky130_fd_sc_hd__a21o_1 _5550_ (.A1(\core_0.decode.oc_alu_mode[2] ),
    .A2(_1571_),
    .B1(\core_0.decode.oc_alu_mode[7] ),
    .X(_2357_));
 sky130_fd_sc_hd__a22o_1 _5551_ (.A1(_1571_),
    .A2(_1776_),
    .B1(_2357_),
    .B2(_1902_),
    .X(_2358_));
 sky130_fd_sc_hd__a221o_1 _5552_ (.A1(_0956_),
    .A2(_1866_),
    .B1(_1949_),
    .B2(\core_0.decode.oc_alu_mode[6] ),
    .C1(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__a41o_1 _5553_ (.A1(_1751_),
    .A2(_1700_),
    .A3(_2097_),
    .A4(_2102_),
    .B1(_2359_),
    .X(_2360_));
 sky130_fd_sc_hd__inv_2 _5554_ (.A(_2360_),
    .Y(_2361_));
 sky130_fd_sc_hd__o221a_1 _5555_ (.A1(_2246_),
    .A2(_2354_),
    .B1(_2355_),
    .B2(_2356_),
    .C1(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__o21ai_1 _5556_ (.A1(_1773_),
    .A2(_2351_),
    .B1(_2362_),
    .Y(_2363_));
 sky130_fd_sc_hd__a31o_2 _5557_ (.A1(_0978_),
    .A2(_2348_),
    .A3(_2349_),
    .B1(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__a21o_1 _5558_ (.A1(_2135_),
    .A2(\core_0.execute.alu_mul_div.mul_res[7] ),
    .B1(_0988_),
    .X(_2365_));
 sky130_fd_sc_hd__a21o_1 _5559_ (.A1(_1784_),
    .A2(_2364_),
    .B1(_2365_),
    .X(_2366_));
 sky130_fd_sc_hd__a22o_4 _5560_ (.A1(\core_0.execute.alu_mul_div.div_cur[7] ),
    .A2(_0960_),
    .B1(_2347_),
    .B2(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__clkbuf_4 _5561_ (.A(_2065_),
    .X(_2368_));
 sky130_fd_sc_hd__clkbuf_4 _5562_ (.A(_2067_),
    .X(_2369_));
 sky130_fd_sc_hd__a22o_1 _5563_ (.A1(\core_0.execute.sreg_irq_pc.o_d[7] ),
    .A2(_2368_),
    .B1(_2369_),
    .B2(\core_0.execute.sreg_scratch.o_d[7] ),
    .X(_2370_));
 sky130_fd_sc_hd__a221o_1 _5564_ (.A1(\core_0.execute.sreg_priv_control.o_d[7] ),
    .A2(_1162_),
    .B1(_2075_),
    .B2(\core_0.execute.pc_high_out[7] ),
    .C1(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__a221o_1 _5565_ (.A1(\core_0.execute.pc_high_buff_out[7] ),
    .A2(_2192_),
    .B1(_2193_),
    .B2(net14),
    .C1(_2371_),
    .X(_2372_));
 sky130_fd_sc_hd__a22o_1 _5566_ (.A1(net85),
    .A2(_2310_),
    .B1(_2372_),
    .B2(_2152_),
    .X(_2373_));
 sky130_fd_sc_hd__mux2_1 _5567_ (.A0(\core_0.execute.sreg_irq_pc.o_d[7] ),
    .A1(_2373_),
    .S(_1788_),
    .X(_2374_));
 sky130_fd_sc_hd__or2b_1 _5568_ (.A(_2317_),
    .B_N(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__a21oi_1 _5569_ (.A1(_2304_),
    .A2(_2315_),
    .B1(_2374_),
    .Y(_2376_));
 sky130_fd_sc_hd__nor2_1 _5570_ (.A(_2159_),
    .B(_2376_),
    .Y(_2377_));
 sky130_fd_sc_hd__a22o_1 _5571_ (.A1(_2159_),
    .A2(_2367_),
    .B1(_2375_),
    .B2(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__mux2_1 _5572_ (.A0(_2378_),
    .A1(net207),
    .S(_2089_),
    .X(_2379_));
 sky130_fd_sc_hd__mux2_1 _5573_ (.A0(_2379_),
    .A1(\core_0.ew_data[7] ),
    .S(_2345_),
    .X(_2380_));
 sky130_fd_sc_hd__clkbuf_1 _5574_ (.A(_2380_),
    .X(_0236_));
 sky130_fd_sc_hd__a21bo_1 _5575_ (.A1(\core_0.execute.alu_mul_div.div_res[8] ),
    .A2(_1696_),
    .B1_N(_0741_),
    .X(_2381_));
 sky130_fd_sc_hd__and2_1 _5576_ (.A(_1901_),
    .B(_1908_),
    .X(_2382_));
 sky130_fd_sc_hd__nor2_1 _5577_ (.A(_1901_),
    .B(_1908_),
    .Y(_2383_));
 sky130_fd_sc_hd__nor4_1 _5578_ (.A(_1865_),
    .B(_1905_),
    .C(_1951_),
    .D(_1956_),
    .Y(_2384_));
 sky130_fd_sc_hd__or2_1 _5579_ (.A(_1773_),
    .B(_1957_),
    .X(_2385_));
 sky130_fd_sc_hd__and2_2 _5580_ (.A(\core_0.decode.oc_alu_mode[3] ),
    .B(_1571_),
    .X(_2386_));
 sky130_fd_sc_hd__a221o_1 _5581_ (.A1(_0934_),
    .A2(_1391_),
    .B1(_1579_),
    .B2(_1775_),
    .C1(_2386_),
    .X(_2387_));
 sky130_fd_sc_hd__a221o_1 _5582_ (.A1(_0998_),
    .A2(_1903_),
    .B1(_1904_),
    .B2(\core_0.decode.oc_alu_mode[9] ),
    .C1(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__a21o_1 _5583_ (.A1(_0928_),
    .A2(_1905_),
    .B1(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__and4_1 _5584_ (.A(_1751_),
    .B(_1700_),
    .C(_1707_),
    .D(_1723_),
    .X(_2390_));
 sky130_fd_sc_hd__a211oi_1 _5585_ (.A1(_1371_),
    .A2(_1762_),
    .B1(_2389_),
    .C1(_2390_),
    .Y(_2391_));
 sky130_fd_sc_hd__o221a_1 _5586_ (.A1(_1986_),
    .A2(_2246_),
    .B1(_2384_),
    .B2(_2385_),
    .C1(_2391_),
    .X(_2392_));
 sky130_fd_sc_hd__o31a_1 _5587_ (.A1(_1774_),
    .A2(_2382_),
    .A3(_2383_),
    .B1(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__nor2_1 _5588_ (.A(_2135_),
    .B(_2393_),
    .Y(_2394_));
 sky130_fd_sc_hd__a211o_1 _5589_ (.A1(_2135_),
    .A2(\core_0.execute.alu_mul_div.mul_res[8] ),
    .B1(_2394_),
    .C1(_0989_),
    .X(_2395_));
 sky130_fd_sc_hd__a22o_4 _5590_ (.A1(\core_0.execute.alu_mul_div.div_cur[8] ),
    .A2(\core_0.execute.alu_mul_div.i_mod ),
    .B1(_2381_),
    .B2(_2395_),
    .X(_2396_));
 sky130_fd_sc_hd__a22o_1 _5591_ (.A1(\core_0.execute.sreg_irq_pc.o_d[8] ),
    .A2(_2368_),
    .B1(_2369_),
    .B2(\core_0.execute.sreg_scratch.o_d[8] ),
    .X(_2397_));
 sky130_fd_sc_hd__a221o_1 _5592_ (.A1(\core_0.execute.sreg_priv_control.o_d[8] ),
    .A2(_1162_),
    .B1(_2076_),
    .B2(net15),
    .C1(_2397_),
    .X(_2398_));
 sky130_fd_sc_hd__a22o_1 _5593_ (.A1(net86),
    .A2(_2310_),
    .B1(_2398_),
    .B2(_2152_),
    .X(_2399_));
 sky130_fd_sc_hd__mux2_1 _5594_ (.A0(\core_0.execute.sreg_irq_pc.o_d[8] ),
    .A1(_2399_),
    .S(_1788_),
    .X(_2400_));
 sky130_fd_sc_hd__xnor2_1 _5595_ (.A(_2375_),
    .B(_2400_),
    .Y(_2401_));
 sky130_fd_sc_hd__mux2_1 _5596_ (.A0(_2396_),
    .A1(_2401_),
    .S(_2087_),
    .X(_2402_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(_2402_),
    .A1(net208),
    .S(_2089_),
    .X(_2403_));
 sky130_fd_sc_hd__mux2_1 _5598_ (.A0(_2403_),
    .A1(\core_0.ew_data[8] ),
    .S(_2345_),
    .X(_2404_));
 sky130_fd_sc_hd__clkbuf_1 _5599_ (.A(_2404_),
    .X(_0237_));
 sky130_fd_sc_hd__inv_2 _5600_ (.A(\core_0.ew_data[9] ),
    .Y(_2405_));
 sky130_fd_sc_hd__a21bo_1 _5601_ (.A1(\core_0.execute.alu_mul_div.div_res[9] ),
    .A2(_1697_),
    .B1_N(_1411_),
    .X(_2406_));
 sky130_fd_sc_hd__nand2_1 _5602_ (.A(_2006_),
    .B(_2281_),
    .Y(_2407_));
 sky130_fd_sc_hd__mux2_1 _5603_ (.A0(_1968_),
    .A1(_1971_),
    .S(_1423_),
    .X(_2408_));
 sky130_fd_sc_hd__mux2_1 _5604_ (.A0(_1972_),
    .A1(_1995_),
    .S(_1423_),
    .X(_2409_));
 sky130_fd_sc_hd__mux2_1 _5605_ (.A0(_2408_),
    .A1(_2409_),
    .S(_1975_),
    .X(_2410_));
 sky130_fd_sc_hd__nand2_1 _5606_ (.A(_1988_),
    .B(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__nor2_1 _5607_ (.A(_1967_),
    .B(_2006_),
    .Y(_2412_));
 sky130_fd_sc_hd__and2b_1 _5608_ (.A_N(_2094_),
    .B(_2412_),
    .X(_2413_));
 sky130_fd_sc_hd__a31o_1 _5609_ (.A1(_1967_),
    .A2(_2407_),
    .A3(_2411_),
    .B1(_2413_),
    .X(_2414_));
 sky130_fd_sc_hd__nor2_1 _5610_ (.A(_2131_),
    .B(_2109_),
    .Y(_2415_));
 sky130_fd_sc_hd__a221o_1 _5611_ (.A1(_0934_),
    .A2(_1482_),
    .B1(_1550_),
    .B2(_1775_),
    .C1(_2386_),
    .X(_2416_));
 sky130_fd_sc_hd__a221o_1 _5612_ (.A1(_0956_),
    .A2(_1858_),
    .B1(_1958_),
    .B2(_0998_),
    .C1(_2416_),
    .X(_2417_));
 sky130_fd_sc_hd__a211o_1 _5613_ (.A1(_0928_),
    .A2(_1860_),
    .B1(_2415_),
    .C1(_2417_),
    .X(_2418_));
 sky130_fd_sc_hd__a21oi_2 _5614_ (.A1(_1707_),
    .A2(_2414_),
    .B1(_2418_),
    .Y(_2419_));
 sky130_fd_sc_hd__o21ai_1 _5615_ (.A1(_1907_),
    .A2(_2382_),
    .B1(_1864_),
    .Y(_2420_));
 sky130_fd_sc_hd__o31a_1 _5616_ (.A1(_1864_),
    .A2(_1907_),
    .A3(_2382_),
    .B1(\core_0.decode.oc_alu_mode[11] ),
    .X(_2421_));
 sky130_fd_sc_hd__o21ai_1 _5617_ (.A1(_1903_),
    .A2(_1957_),
    .B1(_1860_),
    .Y(_2422_));
 sky130_fd_sc_hd__o31a_1 _5618_ (.A1(_1860_),
    .A2(_1903_),
    .A3(_1957_),
    .B1(_0962_),
    .X(_2423_));
 sky130_fd_sc_hd__a22oi_2 _5619_ (.A1(_2420_),
    .A2(_2421_),
    .B1(_2422_),
    .B2(_2423_),
    .Y(_2424_));
 sky130_fd_sc_hd__a21oi_1 _5620_ (.A1(_2419_),
    .A2(_2424_),
    .B1(_0955_),
    .Y(_2425_));
 sky130_fd_sc_hd__a211o_1 _5621_ (.A1(_0955_),
    .A2(\core_0.execute.alu_mul_div.mul_res[9] ),
    .B1(_2425_),
    .C1(_0989_),
    .X(_2426_));
 sky130_fd_sc_hd__a22o_4 _5622_ (.A1(\core_0.execute.alu_mul_div.div_cur[9] ),
    .A2(_0960_),
    .B1(_2406_),
    .B2(_2426_),
    .X(_2427_));
 sky130_fd_sc_hd__nand2_1 _5623_ (.A(_2159_),
    .B(_2427_),
    .Y(_2428_));
 sky130_fd_sc_hd__and2b_1 _5624_ (.A_N(_2375_),
    .B(_2400_),
    .X(_2429_));
 sky130_fd_sc_hd__a22o_1 _5625_ (.A1(\core_0.execute.sreg_irq_pc.o_d[9] ),
    .A2(_2368_),
    .B1(_2369_),
    .B2(\core_0.execute.sreg_scratch.o_d[9] ),
    .X(_2430_));
 sky130_fd_sc_hd__a221o_1 _5626_ (.A1(\core_0.execute.sreg_priv_control.o_d[9] ),
    .A2(_1162_),
    .B1(_2076_),
    .B2(net16),
    .C1(_2430_),
    .X(_2431_));
 sky130_fd_sc_hd__a22o_1 _5627_ (.A1(net87),
    .A2(_2310_),
    .B1(_2431_),
    .B2(_2152_),
    .X(_2432_));
 sky130_fd_sc_hd__and2_1 _5628_ (.A(\core_0.execute.sreg_irq_pc.o_d[9] ),
    .B(\core_0.dec_sreg_irt ),
    .X(_2433_));
 sky130_fd_sc_hd__a21oi_1 _5629_ (.A1(_1789_),
    .A2(_2432_),
    .B1(_2433_),
    .Y(_2434_));
 sky130_fd_sc_hd__xnor2_1 _5630_ (.A(_2429_),
    .B(_2434_),
    .Y(_2435_));
 sky130_fd_sc_hd__a21oi_1 _5631_ (.A1(_2087_),
    .A2(_2435_),
    .B1(_1146_),
    .Y(_2436_));
 sky130_fd_sc_hd__a221o_1 _5632_ (.A1(_1146_),
    .A2(_0598_),
    .B1(_2428_),
    .B2(_2436_),
    .C1(_1836_),
    .X(_2437_));
 sky130_fd_sc_hd__o21ai_1 _5633_ (.A1(_2405_),
    .A2(_0228_),
    .B1(_2437_),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _5634_ (.A(\core_0.ew_data[10] ),
    .Y(_2438_));
 sky130_fd_sc_hd__a21bo_1 _5635_ (.A1(\core_0.execute.alu_mul_div.div_res[10] ),
    .A2(_1697_),
    .B1_N(_1411_),
    .X(_2439_));
 sky130_fd_sc_hd__inv_2 _5636_ (.A(_1926_),
    .Y(_2440_));
 sky130_fd_sc_hd__a21oi_1 _5637_ (.A1(_1911_),
    .A2(_2440_),
    .B1(_1774_),
    .Y(_2441_));
 sky130_fd_sc_hd__o21a_1 _5638_ (.A1(_1911_),
    .A2(_2440_),
    .B1(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__o21a_1 _5639_ (.A1(_1957_),
    .A2(_1959_),
    .B1(_1858_),
    .X(_2443_));
 sky130_fd_sc_hd__nor2_1 _5640_ (.A(_1773_),
    .B(_1960_),
    .Y(_2444_));
 sky130_fd_sc_hd__o21a_1 _5641_ (.A1(_1923_),
    .A2(_2443_),
    .B1(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__a221o_1 _5642_ (.A1(_0934_),
    .A2(_1344_),
    .B1(_1922_),
    .B2(_0956_),
    .C1(_2386_),
    .X(_2446_));
 sky130_fd_sc_hd__nor2_1 _5643_ (.A(_2131_),
    .B(_2175_),
    .Y(_2447_));
 sky130_fd_sc_hd__a221o_1 _5644_ (.A1(_1558_),
    .A2(_1775_),
    .B1(_1921_),
    .B2(_0998_),
    .C1(_2447_),
    .X(_2448_));
 sky130_fd_sc_hd__a211o_1 _5645_ (.A1(_0928_),
    .A2(_1923_),
    .B1(_2446_),
    .C1(_2448_),
    .X(_2449_));
 sky130_fd_sc_hd__and2b_1 _5646_ (.A_N(_2162_),
    .B(_2412_),
    .X(_2450_));
 sky130_fd_sc_hd__inv_2 _5647_ (.A(_1973_),
    .Y(_2451_));
 sky130_fd_sc_hd__mux2_1 _5648_ (.A0(_2451_),
    .A1(_1997_),
    .S(_1975_),
    .X(_2452_));
 sky130_fd_sc_hd__nand2_1 _5649_ (.A(_2006_),
    .B(_2324_),
    .Y(_2453_));
 sky130_fd_sc_hd__o211a_1 _5650_ (.A1(_2006_),
    .A2(_2452_),
    .B1(_2453_),
    .C1(_1967_),
    .X(_2454_));
 sky130_fd_sc_hd__o21a_1 _5651_ (.A1(_2450_),
    .A2(_2454_),
    .B1(_1707_),
    .X(_2455_));
 sky130_fd_sc_hd__or4_4 _5652_ (.A(_2442_),
    .B(_2445_),
    .C(_2449_),
    .D(_2455_),
    .X(_2456_));
 sky130_fd_sc_hd__a21o_1 _5653_ (.A1(_2135_),
    .A2(\core_0.execute.alu_mul_div.mul_res[10] ),
    .B1(_0989_),
    .X(_2457_));
 sky130_fd_sc_hd__a21o_1 _5654_ (.A1(_1784_),
    .A2(_2456_),
    .B1(_2457_),
    .X(_2458_));
 sky130_fd_sc_hd__a22o_4 _5655_ (.A1(\core_0.execute.alu_mul_div.div_cur[10] ),
    .A2(_0960_),
    .B1(_2439_),
    .B2(_2458_),
    .X(_2459_));
 sky130_fd_sc_hd__and2b_1 _5656_ (.A_N(_2434_),
    .B(_2429_),
    .X(_2460_));
 sky130_fd_sc_hd__a22o_1 _5657_ (.A1(\core_0.execute.sreg_irq_pc.o_d[10] ),
    .A2(_2368_),
    .B1(_2369_),
    .B2(\core_0.execute.sreg_scratch.o_d[10] ),
    .X(_2461_));
 sky130_fd_sc_hd__a221o_1 _5658_ (.A1(\core_0.execute.sreg_priv_control.o_d[10] ),
    .A2(_1162_),
    .B1(_2076_),
    .B2(net2),
    .C1(_2461_),
    .X(_2462_));
 sky130_fd_sc_hd__a22o_1 _5659_ (.A1(net73),
    .A2(_2310_),
    .B1(_2462_),
    .B2(_2152_),
    .X(_2463_));
 sky130_fd_sc_hd__nand2_1 _5660_ (.A(\core_0.execute.sreg_irq_pc.o_d[10] ),
    .B(_1038_),
    .Y(_2464_));
 sky130_fd_sc_hd__a21bo_1 _5661_ (.A1(_1789_),
    .A2(_2463_),
    .B1_N(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__nand2_1 _5662_ (.A(_2460_),
    .B(_2465_),
    .Y(_2466_));
 sky130_fd_sc_hd__o21a_1 _5663_ (.A1(_2460_),
    .A2(_2465_),
    .B1(_2087_),
    .X(_2467_));
 sky130_fd_sc_hd__a221oi_2 _5664_ (.A1(_2159_),
    .A2(_2459_),
    .B1(_2466_),
    .B2(_2467_),
    .C1(_1146_),
    .Y(_2468_));
 sky130_fd_sc_hd__a211o_1 _5665_ (.A1(_1146_),
    .A2(_0592_),
    .B1(_1836_),
    .C1(_2468_),
    .X(_2469_));
 sky130_fd_sc_hd__o21ai_1 _5666_ (.A1(_2438_),
    .A2(_0228_),
    .B1(_2469_),
    .Y(_0239_));
 sky130_fd_sc_hd__a21boi_1 _5667_ (.A1(\core_0.execute.alu_mul_div.div_res[11] ),
    .A2(_1696_),
    .B1_N(_0741_),
    .Y(_2470_));
 sky130_fd_sc_hd__a21o_1 _5668_ (.A1(_1911_),
    .A2(_2440_),
    .B1(_1925_),
    .X(_2471_));
 sky130_fd_sc_hd__xnor2_1 _5669_ (.A(_1919_),
    .B(_2471_),
    .Y(_2472_));
 sky130_fd_sc_hd__or3_1 _5670_ (.A(_1916_),
    .B(_1921_),
    .C(_1960_),
    .X(_2473_));
 sky130_fd_sc_hd__o21ai_1 _5671_ (.A1(_1921_),
    .A2(_1960_),
    .B1(_1916_),
    .Y(_2474_));
 sky130_fd_sc_hd__mux2_1 _5672_ (.A0(_1972_),
    .A1(_1995_),
    .S(_1423_),
    .X(_2475_));
 sky130_fd_sc_hd__nor2_1 _5673_ (.A(_0984_),
    .B(_1594_),
    .Y(_2476_));
 sky130_fd_sc_hd__o31a_1 _5674_ (.A1(_1719_),
    .A2(_1721_),
    .A3(_2476_),
    .B1(_1422_),
    .X(_2477_));
 sky130_fd_sc_hd__nor2_1 _5675_ (.A(_0984_),
    .B(_1558_),
    .Y(_2478_));
 sky130_fd_sc_hd__o31a_1 _5676_ (.A1(_1719_),
    .A2(_1721_),
    .A3(_2478_),
    .B1(_1764_),
    .X(_2479_));
 sky130_fd_sc_hd__or3_1 _5677_ (.A(_1981_),
    .B(_2477_),
    .C(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__o211ai_1 _5678_ (.A1(_1975_),
    .A2(_2475_),
    .B1(_2480_),
    .C1(_1988_),
    .Y(_2481_));
 sky130_fd_sc_hd__nand2_1 _5679_ (.A(_2006_),
    .B(_2353_),
    .Y(_2482_));
 sky130_fd_sc_hd__inv_2 _5680_ (.A(_2352_),
    .Y(_2483_));
 sky130_fd_sc_hd__a32o_1 _5681_ (.A1(_1967_),
    .A2(_2481_),
    .A3(_2482_),
    .B1(_2483_),
    .B2(_2412_),
    .X(_2484_));
 sky130_fd_sc_hd__a22o_1 _5682_ (.A1(_1431_),
    .A2(_2217_),
    .B1(_2247_),
    .B2(_2102_),
    .X(_2485_));
 sky130_fd_sc_hd__a221o_1 _5683_ (.A1(_0934_),
    .A2(_1493_),
    .B1(_1594_),
    .B2(_1775_),
    .C1(_2386_),
    .X(_2486_));
 sky130_fd_sc_hd__a221o_1 _5684_ (.A1(_0956_),
    .A2(_1912_),
    .B1(_1915_),
    .B2(_0998_),
    .C1(_2486_),
    .X(_2487_));
 sky130_fd_sc_hd__a221o_1 _5685_ (.A1(_0928_),
    .A2(_1916_),
    .B1(_2485_),
    .B2(_1754_),
    .C1(_2487_),
    .X(_2488_));
 sky130_fd_sc_hd__a21o_1 _5686_ (.A1(_1707_),
    .A2(_2484_),
    .B1(_2488_),
    .X(_2489_));
 sky130_fd_sc_hd__a31o_1 _5687_ (.A1(_0962_),
    .A2(_2473_),
    .A3(_2474_),
    .B1(_2489_),
    .X(_2490_));
 sky130_fd_sc_hd__a21o_1 _5688_ (.A1(_0978_),
    .A2(_2472_),
    .B1(_2490_),
    .X(_2491_));
 sky130_fd_sc_hd__a21o_1 _5689_ (.A1(\core_0.execute.alu_mul_div.i_mul ),
    .A2(\core_0.execute.alu_mul_div.mul_res[11] ),
    .B1(_0988_),
    .X(_2492_));
 sky130_fd_sc_hd__a21oi_1 _5690_ (.A1(_1784_),
    .A2(_2491_),
    .B1(_2492_),
    .Y(_2493_));
 sky130_fd_sc_hd__o2bb2a_2 _5691_ (.A1_N(\core_0.execute.alu_mul_div.div_cur[11] ),
    .A2_N(\core_0.execute.alu_mul_div.i_mod ),
    .B1(_2470_),
    .B2(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__inv_2 _5692_ (.A(_2494_),
    .Y(_2495_));
 sky130_fd_sc_hd__a22o_1 _5693_ (.A1(\core_0.execute.sreg_irq_pc.o_d[11] ),
    .A2(_2368_),
    .B1(_2369_),
    .B2(\core_0.execute.sreg_scratch.o_d[11] ),
    .X(_2496_));
 sky130_fd_sc_hd__a221o_1 _5694_ (.A1(\core_0.execute.sreg_priv_control.o_d[11] ),
    .A2(_1162_),
    .B1(_2076_),
    .B2(net3),
    .C1(_2496_),
    .X(_2497_));
 sky130_fd_sc_hd__a22o_1 _5695_ (.A1(net74),
    .A2(_2310_),
    .B1(_2497_),
    .B2(_2152_),
    .X(_2498_));
 sky130_fd_sc_hd__nand2_1 _5696_ (.A(\core_0.execute.sreg_irq_pc.o_d[11] ),
    .B(_1038_),
    .Y(_2499_));
 sky130_fd_sc_hd__a21bo_1 _5697_ (.A1(_1789_),
    .A2(_2498_),
    .B1_N(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__xnor2_1 _5698_ (.A(_2466_),
    .B(_2500_),
    .Y(_2501_));
 sky130_fd_sc_hd__mux2_1 _5699_ (.A0(_2495_),
    .A1(_2501_),
    .S(_2087_),
    .X(_2502_));
 sky130_fd_sc_hd__mux2_1 _5700_ (.A0(_2502_),
    .A1(net196),
    .S(_2089_),
    .X(_2503_));
 sky130_fd_sc_hd__mux2_1 _5701_ (.A0(_2503_),
    .A1(\core_0.ew_data[11] ),
    .S(_2345_),
    .X(_2504_));
 sky130_fd_sc_hd__clkbuf_1 _5702_ (.A(_2504_),
    .X(_0240_));
 sky130_fd_sc_hd__inv_2 _5703_ (.A(\core_0.ew_data[12] ),
    .Y(_2505_));
 sky130_fd_sc_hd__a21bo_1 _5704_ (.A1(\core_0.execute.alu_mul_div.div_res[12] ),
    .A2(_1697_),
    .B1_N(_1411_),
    .X(_2506_));
 sky130_fd_sc_hd__xor2_1 _5705_ (.A(_1857_),
    .B(_1929_),
    .X(_2507_));
 sky130_fd_sc_hd__and2_1 _5706_ (.A(_1912_),
    .B(_1941_),
    .X(_2508_));
 sky130_fd_sc_hd__a211o_1 _5707_ (.A1(_1916_),
    .A2(_1960_),
    .B1(_2508_),
    .C1(_1854_),
    .X(_2509_));
 sky130_fd_sc_hd__and3b_1 _5708_ (.A_N(_1961_),
    .B(_2509_),
    .C(_0962_),
    .X(_2510_));
 sky130_fd_sc_hd__and2_1 _5709_ (.A(_1707_),
    .B(_2095_),
    .X(_2511_));
 sky130_fd_sc_hd__and2b_1 _5710_ (.A_N(_2248_),
    .B(_2511_),
    .X(_2512_));
 sky130_fd_sc_hd__nor2_1 _5711_ (.A(_2131_),
    .B(_2257_),
    .Y(_2513_));
 sky130_fd_sc_hd__a221o_1 _5712_ (.A1(_0934_),
    .A2(_1400_),
    .B1(_1588_),
    .B2(_1775_),
    .C1(_2386_),
    .X(_2514_));
 sky130_fd_sc_hd__a221o_1 _5713_ (.A1(_0998_),
    .A2(_1852_),
    .B1(_1853_),
    .B2(_0956_),
    .C1(_2514_),
    .X(_2515_));
 sky130_fd_sc_hd__a211o_1 _5714_ (.A1(_0928_),
    .A2(_1854_),
    .B1(_2513_),
    .C1(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__nor2_1 _5715_ (.A(_2006_),
    .B(_1999_),
    .Y(_2517_));
 sky130_fd_sc_hd__a211o_1 _5716_ (.A1(_2006_),
    .A2(_1976_),
    .B1(_2246_),
    .C1(_2517_),
    .X(_2518_));
 sky130_fd_sc_hd__or4b_1 _5717_ (.A(_2510_),
    .B(_2512_),
    .C(_2516_),
    .D_N(_2518_),
    .X(_2519_));
 sky130_fd_sc_hd__a21oi_1 _5718_ (.A1(_0978_),
    .A2(_2507_),
    .B1(_2519_),
    .Y(_2520_));
 sky130_fd_sc_hd__nor2_1 _5719_ (.A(_0955_),
    .B(_2520_),
    .Y(_2521_));
 sky130_fd_sc_hd__a211o_1 _5720_ (.A1(_0955_),
    .A2(\core_0.execute.alu_mul_div.mul_res[12] ),
    .B1(_2521_),
    .C1(_0989_),
    .X(_2522_));
 sky130_fd_sc_hd__a22o_4 _5721_ (.A1(\core_0.execute.alu_mul_div.div_cur[12] ),
    .A2(_0960_),
    .B1(_2506_),
    .B2(_2522_),
    .X(_2523_));
 sky130_fd_sc_hd__nand2_1 _5722_ (.A(_2159_),
    .B(_2523_),
    .Y(_2524_));
 sky130_fd_sc_hd__and3_1 _5723_ (.A(_2460_),
    .B(_2465_),
    .C(_2500_),
    .X(_2525_));
 sky130_fd_sc_hd__a22o_1 _5724_ (.A1(\core_0.execute.sreg_irq_pc.o_d[12] ),
    .A2(_2368_),
    .B1(_2369_),
    .B2(\core_0.execute.sreg_scratch.o_d[12] ),
    .X(_2526_));
 sky130_fd_sc_hd__a221o_1 _5725_ (.A1(\core_0.execute.sreg_priv_control.o_d[12] ),
    .A2(_1162_),
    .B1(_2076_),
    .B2(net4),
    .C1(_2526_),
    .X(_2527_));
 sky130_fd_sc_hd__a22o_1 _5726_ (.A1(net75),
    .A2(_2310_),
    .B1(_2527_),
    .B2(_2152_),
    .X(_2528_));
 sky130_fd_sc_hd__and2_1 _5727_ (.A(\core_0.execute.sreg_irq_pc.o_d[12] ),
    .B(_1038_),
    .X(_2529_));
 sky130_fd_sc_hd__a21oi_1 _5728_ (.A1(_1789_),
    .A2(_2528_),
    .B1(_2529_),
    .Y(_2530_));
 sky130_fd_sc_hd__xnor2_1 _5729_ (.A(_2525_),
    .B(_2530_),
    .Y(_2531_));
 sky130_fd_sc_hd__a21oi_1 _5730_ (.A1(_2087_),
    .A2(_2531_),
    .B1(_1146_),
    .Y(_2532_));
 sky130_fd_sc_hd__a221o_1 _5731_ (.A1(_1146_),
    .A2(_0579_),
    .B1(_2524_),
    .B2(_2532_),
    .C1(_1836_),
    .X(_2533_));
 sky130_fd_sc_hd__o21ai_1 _5732_ (.A1(_2505_),
    .A2(_0228_),
    .B1(_2533_),
    .Y(_0241_));
 sky130_fd_sc_hd__and2b_1 _5733_ (.A_N(_2530_),
    .B(_2525_),
    .X(_2534_));
 sky130_fd_sc_hd__and3_1 _5734_ (.A(net185),
    .B(_1159_),
    .C(_2062_),
    .X(_2535_));
 sky130_fd_sc_hd__a221o_1 _5735_ (.A1(\core_0.execute.sreg_irq_pc.o_d[13] ),
    .A2(_2368_),
    .B1(_2369_),
    .B2(\core_0.execute.sreg_scratch.o_d[13] ),
    .C1(_2535_),
    .X(_2536_));
 sky130_fd_sc_hd__a221o_1 _5736_ (.A1(\core_0.execute.sreg_priv_control.o_d[13] ),
    .A2(_1162_),
    .B1(_2193_),
    .B2(net5),
    .C1(_2536_),
    .X(_2537_));
 sky130_fd_sc_hd__a22o_1 _5737_ (.A1(net76),
    .A2(_2310_),
    .B1(_2537_),
    .B2(_2152_),
    .X(_2538_));
 sky130_fd_sc_hd__mux2_1 _5738_ (.A0(\core_0.execute.sreg_irq_pc.o_d[13] ),
    .A1(_2538_),
    .S(_1789_),
    .X(_2539_));
 sky130_fd_sc_hd__nand2_1 _5739_ (.A(_2534_),
    .B(_2539_),
    .Y(_2540_));
 sky130_fd_sc_hd__o21a_1 _5740_ (.A1(_2534_),
    .A2(_2539_),
    .B1(_2086_),
    .X(_2541_));
 sky130_fd_sc_hd__a21boi_1 _5741_ (.A1(\core_0.execute.alu_mul_div.div_res[13] ),
    .A2(_1697_),
    .B1_N(_1411_),
    .Y(_2542_));
 sky130_fd_sc_hd__a21oi_1 _5742_ (.A1(_1857_),
    .A2(_1929_),
    .B1(_1856_),
    .Y(_2543_));
 sky130_fd_sc_hd__xnor2_2 _5743_ (.A(_1851_),
    .B(_2543_),
    .Y(_2544_));
 sky130_fd_sc_hd__o21ai_1 _5744_ (.A1(_1852_),
    .A2(_1961_),
    .B1(_1848_),
    .Y(_2545_));
 sky130_fd_sc_hd__or3_1 _5745_ (.A(_1848_),
    .B(_1852_),
    .C(_1961_),
    .X(_2546_));
 sky130_fd_sc_hd__and3_1 _5746_ (.A(_0962_),
    .B(_2545_),
    .C(_2546_),
    .X(_2547_));
 sky130_fd_sc_hd__mux2_1 _5747_ (.A0(_1989_),
    .A1(_1992_),
    .S(_2002_),
    .X(_2548_));
 sky130_fd_sc_hd__mux2_1 _5748_ (.A0(_1990_),
    .A1(_2001_),
    .S(_1423_),
    .X(_2549_));
 sky130_fd_sc_hd__mux2_1 _5749_ (.A0(_2548_),
    .A1(_2549_),
    .S(_1975_),
    .X(_2550_));
 sky130_fd_sc_hd__nand2_1 _5750_ (.A(_2006_),
    .B(_2410_),
    .Y(_2551_));
 sky130_fd_sc_hd__o21a_1 _5751_ (.A1(_2006_),
    .A2(_2550_),
    .B1(_2551_),
    .X(_2552_));
 sky130_fd_sc_hd__and2b_1 _5752_ (.A_N(_2282_),
    .B(_2511_),
    .X(_2553_));
 sky130_fd_sc_hd__a221o_1 _5753_ (.A1(_0934_),
    .A2(_1845_),
    .B1(_1601_),
    .B2(_1775_),
    .C1(_2386_),
    .X(_2554_));
 sky130_fd_sc_hd__a221o_1 _5754_ (.A1(_0956_),
    .A2(_1962_),
    .B1(_1847_),
    .B2(_0998_),
    .C1(_2554_),
    .X(_2555_));
 sky130_fd_sc_hd__a21oi_2 _5755_ (.A1(_0928_),
    .A2(_1848_),
    .B1(_2555_),
    .Y(_2556_));
 sky130_fd_sc_hd__o31ai_2 _5756_ (.A1(_1749_),
    .A2(_2131_),
    .A3(_2104_),
    .B1(_2556_),
    .Y(_2557_));
 sky130_fd_sc_hd__a211o_1 _5757_ (.A1(_2321_),
    .A2(_2552_),
    .B1(_2553_),
    .C1(_2557_),
    .X(_2558_));
 sky130_fd_sc_hd__a211oi_4 _5758_ (.A1(_0978_),
    .A2(_2544_),
    .B1(_2547_),
    .C1(_2558_),
    .Y(_2559_));
 sky130_fd_sc_hd__a21oi_1 _5759_ (.A1(_0955_),
    .A2(\core_0.execute.alu_mul_div.mul_res[13] ),
    .B1(_0989_),
    .Y(_2560_));
 sky130_fd_sc_hd__o21a_1 _5760_ (.A1(_0955_),
    .A2(_2559_),
    .B1(_2560_),
    .X(_2561_));
 sky130_fd_sc_hd__o2bb2a_4 _5761_ (.A1_N(\core_0.execute.alu_mul_div.div_cur[13] ),
    .A2_N(_0960_),
    .B1(_2542_),
    .B2(_2561_),
    .X(_2562_));
 sky130_fd_sc_hd__o2bb2a_1 _5762_ (.A1_N(_2540_),
    .A2_N(_2541_),
    .B1(_2087_),
    .B2(_2562_),
    .X(_2563_));
 sky130_fd_sc_hd__nand2_1 _5763_ (.A(_1146_),
    .B(net198),
    .Y(_2564_));
 sky130_fd_sc_hd__o21ai_1 _5764_ (.A1(_1146_),
    .A2(_2563_),
    .B1(_2564_),
    .Y(_2565_));
 sky130_fd_sc_hd__mux2_1 _5765_ (.A0(_2565_),
    .A1(\core_0.ew_data[13] ),
    .S(_2345_),
    .X(_2566_));
 sky130_fd_sc_hd__clkbuf_1 _5766_ (.A(_2566_),
    .X(_0242_));
 sky130_fd_sc_hd__a21o_1 _5767_ (.A1(\core_0.execute.alu_mul_div.div_res[14] ),
    .A2(_0989_),
    .B1(\core_0.execute.alu_mul_div.i_mod ),
    .X(_2567_));
 sky130_fd_sc_hd__and2b_1 _5768_ (.A_N(_1936_),
    .B(_1844_),
    .X(_2568_));
 sky130_fd_sc_hd__nand2_1 _5769_ (.A(_2568_),
    .B(_1931_),
    .Y(_2569_));
 sky130_fd_sc_hd__or2_1 _5770_ (.A(_2568_),
    .B(_1931_),
    .X(_2570_));
 sky130_fd_sc_hd__o21a_1 _5771_ (.A1(_1847_),
    .A2(_1852_),
    .B1(_1962_),
    .X(_2571_));
 sky130_fd_sc_hd__a211o_1 _5772_ (.A1(_1848_),
    .A2(_1961_),
    .B1(_2571_),
    .C1(_1843_),
    .X(_2572_));
 sky130_fd_sc_hd__and3b_1 _5773_ (.A_N(_1963_),
    .B(_2572_),
    .C(_0962_),
    .X(_2573_));
 sky130_fd_sc_hd__mux2_1 _5774_ (.A0(_1991_),
    .A1(_2003_),
    .S(_1975_),
    .X(_2574_));
 sky130_fd_sc_hd__mux2_1 _5775_ (.A0(_2452_),
    .A1(_2574_),
    .S(_1988_),
    .X(_2575_));
 sky130_fd_sc_hd__nor2_1 _5776_ (.A(_2131_),
    .B(_2329_),
    .Y(_2576_));
 sky130_fd_sc_hd__inv_2 _5777_ (.A(_1842_),
    .Y(_2577_));
 sky130_fd_sc_hd__a221o_1 _5778_ (.A1(_0934_),
    .A2(_1331_),
    .B1(_1841_),
    .B2(_1775_),
    .C1(_2386_),
    .X(_2578_));
 sky130_fd_sc_hd__a221o_1 _5779_ (.A1(_0998_),
    .A2(_1840_),
    .B1(_2577_),
    .B2(_0956_),
    .C1(_2578_),
    .X(_2579_));
 sky130_fd_sc_hd__a211o_1 _5780_ (.A1(_0928_),
    .A2(_1843_),
    .B1(_2576_),
    .C1(_2579_),
    .X(_2580_));
 sky130_fd_sc_hd__a221o_1 _5781_ (.A1(_2326_),
    .A2(_2511_),
    .B1(_2575_),
    .B2(_2321_),
    .C1(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__a311o_2 _5782_ (.A1(\core_0.decode.oc_alu_mode[11] ),
    .A2(_2569_),
    .A3(_2570_),
    .B1(_2573_),
    .C1(_2581_),
    .X(_2582_));
 sky130_fd_sc_hd__mux2_1 _5783_ (.A0(\core_0.execute.alu_mul_div.mul_res[14] ),
    .A1(_2582_),
    .S(_1784_),
    .X(_2583_));
 sky130_fd_sc_hd__and2b_1 _5784_ (.A_N(_0989_),
    .B(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__o22a_4 _5785_ (.A1(\core_0.execute.alu_mul_div.div_cur[14] ),
    .A2(_1697_),
    .B1(_2567_),
    .B2(_2584_),
    .X(_2585_));
 sky130_fd_sc_hd__a221o_1 _5786_ (.A1(\core_0.execute.sreg_irq_pc.o_d[14] ),
    .A2(_2368_),
    .B1(_2369_),
    .B2(\core_0.execute.sreg_scratch.o_d[14] ),
    .C1(_2535_),
    .X(_2586_));
 sky130_fd_sc_hd__a221o_1 _5787_ (.A1(\core_0.execute.sreg_priv_control.o_d[14] ),
    .A2(_1162_),
    .B1(_2193_),
    .B2(net6),
    .C1(_2586_),
    .X(_2587_));
 sky130_fd_sc_hd__a22o_1 _5788_ (.A1(net77),
    .A2(_2310_),
    .B1(_2587_),
    .B2(_2152_),
    .X(_2588_));
 sky130_fd_sc_hd__mux2_1 _5789_ (.A0(\core_0.execute.sreg_irq_pc.o_d[14] ),
    .A1(_2588_),
    .S(_1789_),
    .X(_2589_));
 sky130_fd_sc_hd__xnor2_1 _5790_ (.A(_2540_),
    .B(_2589_),
    .Y(_2590_));
 sky130_fd_sc_hd__mux2_1 _5791_ (.A0(_2585_),
    .A1(_2590_),
    .S(_2086_),
    .X(_2591_));
 sky130_fd_sc_hd__mux2_1 _5792_ (.A0(_2591_),
    .A1(net199),
    .S(\core_0.dec_mem_access ),
    .X(_2592_));
 sky130_fd_sc_hd__mux2_1 _5793_ (.A0(_2592_),
    .A1(\core_0.ew_data[14] ),
    .S(_2345_),
    .X(_2593_));
 sky130_fd_sc_hd__clkbuf_1 _5794_ (.A(_2593_),
    .X(_0243_));
 sky130_fd_sc_hd__a21oi_1 _5795_ (.A1(_1844_),
    .A2(_1931_),
    .B1(_1936_),
    .Y(_2594_));
 sky130_fd_sc_hd__nor2_1 _5796_ (.A(_1935_),
    .B(_1938_),
    .Y(_2595_));
 sky130_fd_sc_hd__xnor2_1 _5797_ (.A(_2594_),
    .B(_2595_),
    .Y(_2596_));
 sky130_fd_sc_hd__o21ai_1 _5798_ (.A1(_1840_),
    .A2(_1963_),
    .B1(_1934_),
    .Y(_2597_));
 sky130_fd_sc_hd__o31a_1 _5799_ (.A1(_1934_),
    .A2(_1840_),
    .A3(_1963_),
    .B1(_0962_),
    .X(_2598_));
 sky130_fd_sc_hd__a221o_1 _5800_ (.A1(_0934_),
    .A2(_1839_),
    .B1(_1933_),
    .B2(_0928_),
    .C1(_0956_),
    .X(_2599_));
 sky130_fd_sc_hd__a221o_1 _5801_ (.A1(_0998_),
    .A2(_1940_),
    .B1(_2599_),
    .B2(_1932_),
    .C1(_2386_),
    .X(_2600_));
 sky130_fd_sc_hd__a31o_1 _5802_ (.A1(_1700_),
    .A2(_1754_),
    .A3(_2102_),
    .B1(_2600_),
    .X(_2601_));
 sky130_fd_sc_hd__nand2_1 _5803_ (.A(_1998_),
    .B(_2409_),
    .Y(_2602_));
 sky130_fd_sc_hd__o21a_1 _5804_ (.A1(_1998_),
    .A2(_2548_),
    .B1(_2602_),
    .X(_2603_));
 sky130_fd_sc_hd__nand2_1 _5805_ (.A(_1423_),
    .B(_2004_),
    .Y(_2604_));
 sky130_fd_sc_hd__o21a_1 _5806_ (.A1(_1423_),
    .A2(_2000_),
    .B1(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__mux2_1 _5807_ (.A0(_2549_),
    .A1(_2605_),
    .S(_1975_),
    .X(_2606_));
 sky130_fd_sc_hd__mux2_1 _5808_ (.A0(_2603_),
    .A1(_2606_),
    .S(_1988_),
    .X(_2607_));
 sky130_fd_sc_hd__nand2_1 _5809_ (.A(_2095_),
    .B(_2354_),
    .Y(_2608_));
 sky130_fd_sc_hd__o211a_1 _5810_ (.A1(_2095_),
    .A2(_2607_),
    .B1(_2608_),
    .C1(_1707_),
    .X(_2609_));
 sky130_fd_sc_hd__a211o_1 _5811_ (.A1(_2597_),
    .A2(_2598_),
    .B1(_2601_),
    .C1(_2609_),
    .X(_2610_));
 sky130_fd_sc_hd__a221o_2 _5812_ (.A1(_1542_),
    .A2(_1775_),
    .B1(_2596_),
    .B2(_0978_),
    .C1(_2610_),
    .X(_2611_));
 sky130_fd_sc_hd__a21o_1 _5813_ (.A1(_2135_),
    .A2(\core_0.execute.alu_mul_div.mul_res[15] ),
    .B1(_0988_),
    .X(_2612_));
 sky130_fd_sc_hd__a21o_1 _5814_ (.A1(_1784_),
    .A2(_2611_),
    .B1(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__a21bo_1 _5815_ (.A1(\core_0.execute.alu_mul_div.div_res[15] ),
    .A2(_1696_),
    .B1_N(_0741_),
    .X(_2614_));
 sky130_fd_sc_hd__a22o_4 _5816_ (.A1(\core_0.execute.alu_mul_div.div_cur[15] ),
    .A2(_0960_),
    .B1(_2613_),
    .B2(_2614_),
    .X(_2615_));
 sky130_fd_sc_hd__and3_1 _5817_ (.A(_2534_),
    .B(_2539_),
    .C(_2589_),
    .X(_2616_));
 sky130_fd_sc_hd__a221o_1 _5818_ (.A1(\core_0.execute.sreg_irq_pc.o_d[15] ),
    .A2(_2368_),
    .B1(_2369_),
    .B2(\core_0.execute.sreg_scratch.o_d[15] ),
    .C1(_2535_),
    .X(_2617_));
 sky130_fd_sc_hd__a221o_1 _5819_ (.A1(\core_0.execute.sreg_priv_control.o_d[15] ),
    .A2(_1162_),
    .B1(_2193_),
    .B2(net7),
    .C1(_2617_),
    .X(_2618_));
 sky130_fd_sc_hd__a22o_1 _5820_ (.A1(net78),
    .A2(_2310_),
    .B1(_2618_),
    .B2(_2152_),
    .X(_2619_));
 sky130_fd_sc_hd__mux2_1 _5821_ (.A0(\core_0.execute.sreg_irq_pc.o_d[15] ),
    .A1(_2619_),
    .S(_1789_),
    .X(_2620_));
 sky130_fd_sc_hd__or2_1 _5822_ (.A(_2616_),
    .B(_2620_),
    .X(_2621_));
 sky130_fd_sc_hd__a21oi_1 _5823_ (.A1(_2616_),
    .A2(_2620_),
    .B1(_2159_),
    .Y(_2622_));
 sky130_fd_sc_hd__a22o_1 _5824_ (.A1(_2159_),
    .A2(_2615_),
    .B1(_2621_),
    .B2(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__mux2_1 _5825_ (.A0(_2623_),
    .A1(net200),
    .S(\core_0.dec_mem_access ),
    .X(_2624_));
 sky130_fd_sc_hd__mux2_1 _5826_ (.A0(_2624_),
    .A1(\core_0.ew_data[15] ),
    .S(_2345_),
    .X(_2625_));
 sky130_fd_sc_hd__clkbuf_1 _5827_ (.A(_2625_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5828_ (.A0(_1787_),
    .A1(\core_0.ew_addr[0] ),
    .S(_2345_),
    .X(_2626_));
 sky130_fd_sc_hd__clkbuf_1 _5829_ (.A(_2626_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5830_ (.A0(_2138_),
    .A1(net116),
    .S(_2345_),
    .X(_2627_));
 sky130_fd_sc_hd__clkbuf_1 _5831_ (.A(_2627_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5832_ (.A0(_2187_),
    .A1(net123),
    .S(_2345_),
    .X(_2628_));
 sky130_fd_sc_hd__clkbuf_1 _5833_ (.A(_2628_),
    .X(_0247_));
 sky130_fd_sc_hd__buf_4 _5834_ (.A(_1835_),
    .X(_2629_));
 sky130_fd_sc_hd__mux2_1 _5835_ (.A0(_2241_),
    .A1(net124),
    .S(_2629_),
    .X(_2630_));
 sky130_fd_sc_hd__clkbuf_1 _5836_ (.A(_2630_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _5837_ (.A0(_2266_),
    .A1(net125),
    .S(_2629_),
    .X(_2631_));
 sky130_fd_sc_hd__clkbuf_1 _5838_ (.A(_2631_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _5839_ (.A0(_2298_),
    .A1(net126),
    .S(_2629_),
    .X(_2632_));
 sky130_fd_sc_hd__clkbuf_1 _5840_ (.A(_2632_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5841_ (.A0(_2341_),
    .A1(net127),
    .S(_2629_),
    .X(_2633_));
 sky130_fd_sc_hd__clkbuf_1 _5842_ (.A(_2633_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5843_ (.A0(_2367_),
    .A1(net128),
    .S(_2629_),
    .X(_2634_));
 sky130_fd_sc_hd__clkbuf_1 _5844_ (.A(_2634_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5845_ (.A0(_2396_),
    .A1(net129),
    .S(_2629_),
    .X(_2635_));
 sky130_fd_sc_hd__clkbuf_1 _5846_ (.A(_2635_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5847_ (.A0(_2427_),
    .A1(net130),
    .S(_2629_),
    .X(_2636_));
 sky130_fd_sc_hd__clkbuf_1 _5848_ (.A(_2636_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5849_ (.A0(_2459_),
    .A1(net131),
    .S(_2629_),
    .X(_2637_));
 sky130_fd_sc_hd__clkbuf_1 _5850_ (.A(_2637_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5851_ (.A0(_2495_),
    .A1(net117),
    .S(_2629_),
    .X(_2638_));
 sky130_fd_sc_hd__clkbuf_1 _5852_ (.A(_2638_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5853_ (.A0(_2523_),
    .A1(net118),
    .S(_2629_),
    .X(_2639_));
 sky130_fd_sc_hd__clkbuf_1 _5854_ (.A(_2639_),
    .X(_0257_));
 sky130_fd_sc_hd__nand2_1 _5855_ (.A(net119),
    .B(_1836_),
    .Y(_2640_));
 sky130_fd_sc_hd__o21ai_1 _5856_ (.A1(_1836_),
    .A2(_2562_),
    .B1(_2640_),
    .Y(_0258_));
 sky130_fd_sc_hd__buf_4 _5857_ (.A(_1835_),
    .X(_2641_));
 sky130_fd_sc_hd__mux2_1 _5858_ (.A0(_2585_),
    .A1(net120),
    .S(_2641_),
    .X(_2642_));
 sky130_fd_sc_hd__clkbuf_1 _5859_ (.A(_2642_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5860_ (.A0(_2615_),
    .A1(net121),
    .S(_2641_),
    .X(_2643_));
 sky130_fd_sc_hd__clkbuf_1 _5861_ (.A(_2643_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5862_ (.A0(\core_0.dec_rf_ie[0] ),
    .A1(\core_0.ew_reg_ie[0] ),
    .S(_2641_),
    .X(_2644_));
 sky130_fd_sc_hd__clkbuf_1 _5863_ (.A(_2644_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5864_ (.A0(\core_0.dec_rf_ie[1] ),
    .A1(\core_0.ew_reg_ie[1] ),
    .S(_2641_),
    .X(_2645_));
 sky130_fd_sc_hd__clkbuf_1 _5865_ (.A(_2645_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5866_ (.A0(\core_0.dec_rf_ie[2] ),
    .A1(\core_0.ew_reg_ie[2] ),
    .S(_2641_),
    .X(_2646_));
 sky130_fd_sc_hd__clkbuf_1 _5867_ (.A(_2646_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5868_ (.A0(\core_0.dec_rf_ie[3] ),
    .A1(\core_0.ew_reg_ie[3] ),
    .S(_2641_),
    .X(_2647_));
 sky130_fd_sc_hd__clkbuf_1 _5869_ (.A(_2647_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _5870_ (.A0(\core_0.dec_rf_ie[4] ),
    .A1(\core_0.ew_reg_ie[4] ),
    .S(_2641_),
    .X(_2648_));
 sky130_fd_sc_hd__clkbuf_1 _5871_ (.A(_2648_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5872_ (.A0(\core_0.dec_rf_ie[5] ),
    .A1(\core_0.ew_reg_ie[5] ),
    .S(_2641_),
    .X(_2649_));
 sky130_fd_sc_hd__clkbuf_1 _5873_ (.A(_2649_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _5874_ (.A0(\core_0.dec_rf_ie[6] ),
    .A1(\core_0.ew_reg_ie[6] ),
    .S(_2641_),
    .X(_2650_));
 sky130_fd_sc_hd__clkbuf_1 _5875_ (.A(_2650_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _5876_ (.A0(\core_0.dec_rf_ie[7] ),
    .A1(\core_0.ew_reg_ie[7] ),
    .S(_2641_),
    .X(_2651_));
 sky130_fd_sc_hd__clkbuf_1 _5877_ (.A(_2651_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5878_ (.A0(_1146_),
    .A1(_1318_),
    .S(_1835_),
    .X(_2652_));
 sky130_fd_sc_hd__clkbuf_1 _5879_ (.A(_2652_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5880_ (.A0(\core_0.dec_mem_width ),
    .A1(\core_0.ew_mem_width ),
    .S(_1835_),
    .X(_2653_));
 sky130_fd_sc_hd__clkbuf_1 _5881_ (.A(_2653_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5882_ (.A0(_0721_),
    .A1(net155),
    .S(_1835_),
    .X(_2654_));
 sky130_fd_sc_hd__clkbuf_1 _5883_ (.A(_2654_),
    .X(_0271_));
 sky130_fd_sc_hd__nor2_1 _5884_ (.A(_1128_),
    .B(_1158_),
    .Y(_0272_));
 sky130_fd_sc_hd__mux2_8 _5885_ (.A0(\core_0.ew_submit ),
    .A1(net20),
    .S(\core_0.ew_mem_access ),
    .X(_2655_));
 sky130_fd_sc_hd__buf_8 _5886_ (.A(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__nand2_4 _5887_ (.A(\core_0.ew_reg_ie[7] ),
    .B(_2656_),
    .Y(_2657_));
 sky130_fd_sc_hd__mux2_1 _5888_ (.A0(net35),
    .A1(net21),
    .S(_1006_),
    .X(_2658_));
 sky130_fd_sc_hd__mux2_1 _5889_ (.A0(\core_0.ew_data[0] ),
    .A1(_2658_),
    .S(_1317_),
    .X(_2659_));
 sky130_fd_sc_hd__buf_6 _5890_ (.A(_2659_),
    .X(_2660_));
 sky130_fd_sc_hd__and2_2 _5891_ (.A(\core_0.ew_reg_ie[7] ),
    .B(_2655_),
    .X(_2661_));
 sky130_fd_sc_hd__buf_2 _5892_ (.A(_2661_),
    .X(_2662_));
 sky130_fd_sc_hd__or2_1 _5893_ (.A(\core_0.execute.rf.reg_outputs[7][0] ),
    .B(_2662_),
    .X(_2663_));
 sky130_fd_sc_hd__clkbuf_4 _5894_ (.A(_1314_),
    .X(_2664_));
 sky130_fd_sc_hd__o211a_1 _5895_ (.A1(_2657_),
    .A2(_2660_),
    .B1(_2663_),
    .C1(_2664_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5896_ (.A0(net36),
    .A1(net28),
    .S(_1006_),
    .X(_2665_));
 sky130_fd_sc_hd__mux2_1 _5897_ (.A0(\core_0.ew_data[1] ),
    .A1(_2665_),
    .S(_1317_),
    .X(_2666_));
 sky130_fd_sc_hd__buf_6 _5898_ (.A(_2666_),
    .X(_2667_));
 sky130_fd_sc_hd__or2_1 _5899_ (.A(\core_0.execute.rf.reg_outputs[7][1] ),
    .B(_2662_),
    .X(_2668_));
 sky130_fd_sc_hd__o211a_1 _5900_ (.A1(_2657_),
    .A2(_2667_),
    .B1(_2668_),
    .C1(_2664_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5901_ (.A0(net22),
    .A1(net29),
    .S(_1005_),
    .X(_2669_));
 sky130_fd_sc_hd__mux2_1 _5902_ (.A0(\core_0.ew_data[2] ),
    .A1(_2669_),
    .S(_1317_),
    .X(_2670_));
 sky130_fd_sc_hd__buf_6 _5903_ (.A(_2670_),
    .X(_2671_));
 sky130_fd_sc_hd__or2_1 _5904_ (.A(\core_0.execute.rf.reg_outputs[7][2] ),
    .B(_2662_),
    .X(_2672_));
 sky130_fd_sc_hd__o211a_1 _5905_ (.A1(_2657_),
    .A2(_2671_),
    .B1(_2672_),
    .C1(_2664_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5906_ (.A0(net23),
    .A1(net30),
    .S(_1005_),
    .X(_2673_));
 sky130_fd_sc_hd__mux2_1 _5907_ (.A0(\core_0.ew_data[3] ),
    .A1(_2673_),
    .S(_1317_),
    .X(_2674_));
 sky130_fd_sc_hd__buf_6 _5908_ (.A(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__or2_1 _5909_ (.A(\core_0.execute.rf.reg_outputs[7][3] ),
    .B(_2662_),
    .X(_2676_));
 sky130_fd_sc_hd__o211a_1 _5910_ (.A1(_2657_),
    .A2(_2675_),
    .B1(_2676_),
    .C1(_2664_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5911_ (.A0(net24),
    .A1(net31),
    .S(_1005_),
    .X(_2677_));
 sky130_fd_sc_hd__mux2_1 _5912_ (.A0(\core_0.ew_data[4] ),
    .A1(_2677_),
    .S(_1317_),
    .X(_2678_));
 sky130_fd_sc_hd__buf_6 _5913_ (.A(_2678_),
    .X(_2679_));
 sky130_fd_sc_hd__or2_1 _5914_ (.A(\core_0.execute.rf.reg_outputs[7][4] ),
    .B(_2661_),
    .X(_2680_));
 sky130_fd_sc_hd__o211a_1 _5915_ (.A1(_2657_),
    .A2(_2679_),
    .B1(_2680_),
    .C1(_2664_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5916_ (.A0(net25),
    .A1(net32),
    .S(_1005_),
    .X(_2681_));
 sky130_fd_sc_hd__mux2_1 _5917_ (.A0(\core_0.ew_data[5] ),
    .A1(_2681_),
    .S(_1317_),
    .X(_2682_));
 sky130_fd_sc_hd__buf_6 _5918_ (.A(_2682_),
    .X(_2683_));
 sky130_fd_sc_hd__or2_1 _5919_ (.A(\core_0.execute.rf.reg_outputs[7][5] ),
    .B(_2661_),
    .X(_2684_));
 sky130_fd_sc_hd__o211a_1 _5920_ (.A1(_2657_),
    .A2(_2683_),
    .B1(_2684_),
    .C1(_2664_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5921_ (.A0(net26),
    .A1(net33),
    .S(_1005_),
    .X(_2685_));
 sky130_fd_sc_hd__mux2_1 _5922_ (.A0(\core_0.ew_data[6] ),
    .A1(_2685_),
    .S(_1317_),
    .X(_2686_));
 sky130_fd_sc_hd__buf_6 _5923_ (.A(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__or2_1 _5924_ (.A(\core_0.execute.rf.reg_outputs[7][6] ),
    .B(_2661_),
    .X(_2688_));
 sky130_fd_sc_hd__o211a_1 _5925_ (.A1(_2657_),
    .A2(_2687_),
    .B1(_2688_),
    .C1(_2664_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5926_ (.A0(net27),
    .A1(net34),
    .S(_1005_),
    .X(_2689_));
 sky130_fd_sc_hd__mux2_1 _5927_ (.A0(\core_0.ew_data[7] ),
    .A1(_2689_),
    .S(_1317_),
    .X(_2690_));
 sky130_fd_sc_hd__buf_6 _5928_ (.A(_2690_),
    .X(_2691_));
 sky130_fd_sc_hd__or2_1 _5929_ (.A(\core_0.execute.rf.reg_outputs[7][7] ),
    .B(_2661_),
    .X(_2692_));
 sky130_fd_sc_hd__o211a_1 _5930_ (.A1(_2657_),
    .A2(_2691_),
    .B1(_2692_),
    .C1(_2664_),
    .X(_0280_));
 sky130_fd_sc_hd__buf_2 _5931_ (.A(_2661_),
    .X(_2693_));
 sky130_fd_sc_hd__and2b_1 _5932_ (.A_N(\core_0.ew_mem_width ),
    .B(_1317_),
    .X(_2694_));
 sky130_fd_sc_hd__clkbuf_4 _5933_ (.A(_2694_),
    .X(_2695_));
 sky130_fd_sc_hd__inv_2 _5934_ (.A(\core_0.ew_data[8] ),
    .Y(_2696_));
 sky130_fd_sc_hd__o2bb2a_4 _5935_ (.A1_N(net35),
    .A2_N(_2695_),
    .B1(_2696_),
    .B2(_1318_),
    .X(_2697_));
 sky130_fd_sc_hd__nand2_1 _5936_ (.A(_2693_),
    .B(_2697_),
    .Y(_2698_));
 sky130_fd_sc_hd__o211a_1 _5937_ (.A1(\core_0.execute.rf.reg_outputs[7][8] ),
    .A2(_2693_),
    .B1(_2698_),
    .C1(_2664_),
    .X(_0281_));
 sky130_fd_sc_hd__o2bb2a_4 _5938_ (.A1_N(net36),
    .A2_N(_2695_),
    .B1(_2405_),
    .B2(_1318_),
    .X(_2699_));
 sky130_fd_sc_hd__nand2_1 _5939_ (.A(_2693_),
    .B(_2699_),
    .Y(_2700_));
 sky130_fd_sc_hd__o211a_1 _5940_ (.A1(\core_0.execute.rf.reg_outputs[7][9] ),
    .A2(_2693_),
    .B1(_2700_),
    .C1(_2664_),
    .X(_0282_));
 sky130_fd_sc_hd__o2bb2a_4 _5941_ (.A1_N(net22),
    .A2_N(_2695_),
    .B1(_2438_),
    .B2(_1318_),
    .X(_2701_));
 sky130_fd_sc_hd__nand2_1 _5942_ (.A(_2662_),
    .B(_2701_),
    .Y(_2702_));
 sky130_fd_sc_hd__buf_2 _5943_ (.A(_1314_),
    .X(_2703_));
 sky130_fd_sc_hd__o211a_1 _5944_ (.A1(\core_0.execute.rf.reg_outputs[7][10] ),
    .A2(_2693_),
    .B1(_2702_),
    .C1(_2703_),
    .X(_0283_));
 sky130_fd_sc_hd__inv_2 _5945_ (.A(\core_0.ew_data[11] ),
    .Y(_2704_));
 sky130_fd_sc_hd__o2bb2a_4 _5946_ (.A1_N(net23),
    .A2_N(_2695_),
    .B1(_2704_),
    .B2(_1318_),
    .X(_2705_));
 sky130_fd_sc_hd__nand2_1 _5947_ (.A(_2662_),
    .B(_2705_),
    .Y(_2706_));
 sky130_fd_sc_hd__o211a_1 _5948_ (.A1(\core_0.execute.rf.reg_outputs[7][11] ),
    .A2(_2693_),
    .B1(_2706_),
    .C1(_2703_),
    .X(_0284_));
 sky130_fd_sc_hd__o2bb2a_4 _5949_ (.A1_N(net24),
    .A2_N(_2695_),
    .B1(_2505_),
    .B2(_1318_),
    .X(_2707_));
 sky130_fd_sc_hd__nand2_1 _5950_ (.A(_2662_),
    .B(_2707_),
    .Y(_2708_));
 sky130_fd_sc_hd__o211a_1 _5951_ (.A1(\core_0.execute.rf.reg_outputs[7][12] ),
    .A2(_2693_),
    .B1(_2708_),
    .C1(_2703_),
    .X(_0285_));
 sky130_fd_sc_hd__inv_2 _5952_ (.A(\core_0.ew_data[13] ),
    .Y(_2709_));
 sky130_fd_sc_hd__o2bb2a_4 _5953_ (.A1_N(net25),
    .A2_N(_2695_),
    .B1(_2709_),
    .B2(_1318_),
    .X(_2710_));
 sky130_fd_sc_hd__nand2_1 _5954_ (.A(_2662_),
    .B(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__o211a_1 _5955_ (.A1(\core_0.execute.rf.reg_outputs[7][13] ),
    .A2(_2693_),
    .B1(_2711_),
    .C1(_2703_),
    .X(_0286_));
 sky130_fd_sc_hd__inv_2 _5956_ (.A(\core_0.ew_data[14] ),
    .Y(_2712_));
 sky130_fd_sc_hd__o2bb2a_4 _5957_ (.A1_N(net26),
    .A2_N(_2695_),
    .B1(_2712_),
    .B2(_1318_),
    .X(_2713_));
 sky130_fd_sc_hd__nand2_1 _5958_ (.A(_2662_),
    .B(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__o211a_1 _5959_ (.A1(\core_0.execute.rf.reg_outputs[7][14] ),
    .A2(_2693_),
    .B1(_2714_),
    .C1(_2703_),
    .X(_0287_));
 sky130_fd_sc_hd__inv_2 _5960_ (.A(\core_0.ew_data[15] ),
    .Y(_2715_));
 sky130_fd_sc_hd__o2bb2a_4 _5961_ (.A1_N(net27),
    .A2_N(_2695_),
    .B1(_2715_),
    .B2(_1318_),
    .X(_2716_));
 sky130_fd_sc_hd__nand2_1 _5962_ (.A(_2662_),
    .B(_2716_),
    .Y(_2717_));
 sky130_fd_sc_hd__o211a_1 _5963_ (.A1(\core_0.execute.rf.reg_outputs[7][15] ),
    .A2(_2693_),
    .B1(_2717_),
    .C1(_2703_),
    .X(_0288_));
 sky130_fd_sc_hd__nand2_4 _5964_ (.A(\core_0.ew_reg_ie[6] ),
    .B(_2656_),
    .Y(_2718_));
 sky130_fd_sc_hd__and2_2 _5965_ (.A(\core_0.ew_reg_ie[6] ),
    .B(_2656_),
    .X(_2719_));
 sky130_fd_sc_hd__buf_2 _5966_ (.A(_2719_),
    .X(_2720_));
 sky130_fd_sc_hd__or2_1 _5967_ (.A(\core_0.execute.rf.reg_outputs[6][0] ),
    .B(_2720_),
    .X(_2721_));
 sky130_fd_sc_hd__o211a_1 _5968_ (.A1(_2660_),
    .A2(_2718_),
    .B1(_2721_),
    .C1(_2703_),
    .X(_0289_));
 sky130_fd_sc_hd__or2_1 _5969_ (.A(\core_0.execute.rf.reg_outputs[6][1] ),
    .B(_2720_),
    .X(_2722_));
 sky130_fd_sc_hd__o211a_1 _5970_ (.A1(_2667_),
    .A2(_2718_),
    .B1(_2722_),
    .C1(_2703_),
    .X(_0290_));
 sky130_fd_sc_hd__or2_1 _5971_ (.A(\core_0.execute.rf.reg_outputs[6][2] ),
    .B(_2720_),
    .X(_2723_));
 sky130_fd_sc_hd__o211a_1 _5972_ (.A1(_2671_),
    .A2(_2718_),
    .B1(_2723_),
    .C1(_2703_),
    .X(_0291_));
 sky130_fd_sc_hd__or2_1 _5973_ (.A(\core_0.execute.rf.reg_outputs[6][3] ),
    .B(_2720_),
    .X(_2724_));
 sky130_fd_sc_hd__o211a_1 _5974_ (.A1(_2675_),
    .A2(_2718_),
    .B1(_2724_),
    .C1(_2703_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _5975_ (.A(\core_0.execute.rf.reg_outputs[6][4] ),
    .B(_2719_),
    .X(_2725_));
 sky130_fd_sc_hd__clkbuf_4 _5976_ (.A(_1314_),
    .X(_2726_));
 sky130_fd_sc_hd__o211a_1 _5977_ (.A1(_2679_),
    .A2(_2718_),
    .B1(_2725_),
    .C1(_2726_),
    .X(_0293_));
 sky130_fd_sc_hd__or2_1 _5978_ (.A(\core_0.execute.rf.reg_outputs[6][5] ),
    .B(_2719_),
    .X(_2727_));
 sky130_fd_sc_hd__o211a_1 _5979_ (.A1(_2683_),
    .A2(_2718_),
    .B1(_2727_),
    .C1(_2726_),
    .X(_0294_));
 sky130_fd_sc_hd__or2_1 _5980_ (.A(\core_0.execute.rf.reg_outputs[6][6] ),
    .B(_2719_),
    .X(_2728_));
 sky130_fd_sc_hd__o211a_1 _5981_ (.A1(_2687_),
    .A2(_2718_),
    .B1(_2728_),
    .C1(_2726_),
    .X(_0295_));
 sky130_fd_sc_hd__or2_1 _5982_ (.A(\core_0.execute.rf.reg_outputs[6][7] ),
    .B(_2719_),
    .X(_2729_));
 sky130_fd_sc_hd__o211a_1 _5983_ (.A1(_2691_),
    .A2(_2718_),
    .B1(_2729_),
    .C1(_2726_),
    .X(_0296_));
 sky130_fd_sc_hd__buf_2 _5984_ (.A(_2719_),
    .X(_2730_));
 sky130_fd_sc_hd__nand2_1 _5985_ (.A(_2697_),
    .B(_2730_),
    .Y(_2731_));
 sky130_fd_sc_hd__o211a_1 _5986_ (.A1(\core_0.execute.rf.reg_outputs[6][8] ),
    .A2(_2730_),
    .B1(_2731_),
    .C1(_2726_),
    .X(_0297_));
 sky130_fd_sc_hd__nand2_1 _5987_ (.A(_2699_),
    .B(_2730_),
    .Y(_2732_));
 sky130_fd_sc_hd__o211a_1 _5988_ (.A1(\core_0.execute.rf.reg_outputs[6][9] ),
    .A2(_2730_),
    .B1(_2732_),
    .C1(_2726_),
    .X(_0298_));
 sky130_fd_sc_hd__nand2_1 _5989_ (.A(_2701_),
    .B(_2720_),
    .Y(_2733_));
 sky130_fd_sc_hd__o211a_1 _5990_ (.A1(\core_0.execute.rf.reg_outputs[6][10] ),
    .A2(_2730_),
    .B1(_2733_),
    .C1(_2726_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _5991_ (.A(_2705_),
    .B(_2720_),
    .Y(_2734_));
 sky130_fd_sc_hd__o211a_1 _5992_ (.A1(\core_0.execute.rf.reg_outputs[6][11] ),
    .A2(_2730_),
    .B1(_2734_),
    .C1(_2726_),
    .X(_0300_));
 sky130_fd_sc_hd__nand2_1 _5993_ (.A(_2707_),
    .B(_2720_),
    .Y(_2735_));
 sky130_fd_sc_hd__o211a_1 _5994_ (.A1(\core_0.execute.rf.reg_outputs[6][12] ),
    .A2(_2730_),
    .B1(_2735_),
    .C1(_2726_),
    .X(_0301_));
 sky130_fd_sc_hd__nand2_1 _5995_ (.A(_2710_),
    .B(_2720_),
    .Y(_2736_));
 sky130_fd_sc_hd__o211a_1 _5996_ (.A1(\core_0.execute.rf.reg_outputs[6][13] ),
    .A2(_2730_),
    .B1(_2736_),
    .C1(_2726_),
    .X(_0302_));
 sky130_fd_sc_hd__nand2_1 _5997_ (.A(_2713_),
    .B(_2720_),
    .Y(_2737_));
 sky130_fd_sc_hd__clkbuf_4 _5998_ (.A(_1314_),
    .X(_2738_));
 sky130_fd_sc_hd__o211a_1 _5999_ (.A1(\core_0.execute.rf.reg_outputs[6][14] ),
    .A2(_2730_),
    .B1(_2737_),
    .C1(_2738_),
    .X(_0303_));
 sky130_fd_sc_hd__nand2_1 _6000_ (.A(_2716_),
    .B(_2720_),
    .Y(_2739_));
 sky130_fd_sc_hd__o211a_1 _6001_ (.A1(\core_0.execute.rf.reg_outputs[6][15] ),
    .A2(_2730_),
    .B1(_2739_),
    .C1(_2738_),
    .X(_0304_));
 sky130_fd_sc_hd__nand2_4 _6002_ (.A(\core_0.ew_reg_ie[5] ),
    .B(_2656_),
    .Y(_2740_));
 sky130_fd_sc_hd__and2_2 _6003_ (.A(\core_0.ew_reg_ie[5] ),
    .B(_2656_),
    .X(_2741_));
 sky130_fd_sc_hd__buf_2 _6004_ (.A(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__or2_1 _6005_ (.A(\core_0.execute.rf.reg_outputs[5][0] ),
    .B(_2742_),
    .X(_2743_));
 sky130_fd_sc_hd__o211a_1 _6006_ (.A1(_2660_),
    .A2(_2740_),
    .B1(_2743_),
    .C1(_2738_),
    .X(_0305_));
 sky130_fd_sc_hd__or2_1 _6007_ (.A(\core_0.execute.rf.reg_outputs[5][1] ),
    .B(_2742_),
    .X(_2744_));
 sky130_fd_sc_hd__o211a_1 _6008_ (.A1(_2667_),
    .A2(_2740_),
    .B1(_2744_),
    .C1(_2738_),
    .X(_0306_));
 sky130_fd_sc_hd__or2_1 _6009_ (.A(\core_0.execute.rf.reg_outputs[5][2] ),
    .B(_2742_),
    .X(_2745_));
 sky130_fd_sc_hd__o211a_1 _6010_ (.A1(_2671_),
    .A2(_2740_),
    .B1(_2745_),
    .C1(_2738_),
    .X(_0307_));
 sky130_fd_sc_hd__or2_1 _6011_ (.A(\core_0.execute.rf.reg_outputs[5][3] ),
    .B(_2742_),
    .X(_2746_));
 sky130_fd_sc_hd__o211a_1 _6012_ (.A1(_2675_),
    .A2(_2740_),
    .B1(_2746_),
    .C1(_2738_),
    .X(_0308_));
 sky130_fd_sc_hd__or2_1 _6013_ (.A(\core_0.execute.rf.reg_outputs[5][4] ),
    .B(_2741_),
    .X(_2747_));
 sky130_fd_sc_hd__o211a_1 _6014_ (.A1(_2679_),
    .A2(_2740_),
    .B1(_2747_),
    .C1(_2738_),
    .X(_0309_));
 sky130_fd_sc_hd__or2_1 _6015_ (.A(\core_0.execute.rf.reg_outputs[5][5] ),
    .B(_2741_),
    .X(_2748_));
 sky130_fd_sc_hd__o211a_1 _6016_ (.A1(_2683_),
    .A2(_2740_),
    .B1(_2748_),
    .C1(_2738_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _6017_ (.A(\core_0.execute.rf.reg_outputs[5][6] ),
    .B(_2741_),
    .X(_2749_));
 sky130_fd_sc_hd__o211a_1 _6018_ (.A1(_2687_),
    .A2(_2740_),
    .B1(_2749_),
    .C1(_2738_),
    .X(_0311_));
 sky130_fd_sc_hd__or2_1 _6019_ (.A(\core_0.execute.rf.reg_outputs[5][7] ),
    .B(_2741_),
    .X(_2750_));
 sky130_fd_sc_hd__o211a_1 _6020_ (.A1(_2691_),
    .A2(_2740_),
    .B1(_2750_),
    .C1(_2738_),
    .X(_0312_));
 sky130_fd_sc_hd__buf_2 _6021_ (.A(_2741_),
    .X(_2751_));
 sky130_fd_sc_hd__nand2_1 _6022_ (.A(_2697_),
    .B(_2751_),
    .Y(_2752_));
 sky130_fd_sc_hd__clkbuf_4 _6023_ (.A(_1314_),
    .X(_2753_));
 sky130_fd_sc_hd__o211a_1 _6024_ (.A1(\core_0.execute.rf.reg_outputs[5][8] ),
    .A2(_2751_),
    .B1(_2752_),
    .C1(_2753_),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _6025_ (.A(_2699_),
    .B(_2751_),
    .Y(_2754_));
 sky130_fd_sc_hd__o211a_1 _6026_ (.A1(\core_0.execute.rf.reg_outputs[5][9] ),
    .A2(_2751_),
    .B1(_2754_),
    .C1(_2753_),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _6027_ (.A(_2701_),
    .B(_2742_),
    .Y(_2755_));
 sky130_fd_sc_hd__o211a_1 _6028_ (.A1(\core_0.execute.rf.reg_outputs[5][10] ),
    .A2(_2751_),
    .B1(_2755_),
    .C1(_2753_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_1 _6029_ (.A(_2705_),
    .B(_2742_),
    .Y(_2756_));
 sky130_fd_sc_hd__o211a_1 _6030_ (.A1(\core_0.execute.rf.reg_outputs[5][11] ),
    .A2(_2751_),
    .B1(_2756_),
    .C1(_2753_),
    .X(_0316_));
 sky130_fd_sc_hd__nand2_1 _6031_ (.A(_2707_),
    .B(_2742_),
    .Y(_2757_));
 sky130_fd_sc_hd__o211a_1 _6032_ (.A1(\core_0.execute.rf.reg_outputs[5][12] ),
    .A2(_2751_),
    .B1(_2757_),
    .C1(_2753_),
    .X(_0317_));
 sky130_fd_sc_hd__nand2_1 _6033_ (.A(_2710_),
    .B(_2742_),
    .Y(_2758_));
 sky130_fd_sc_hd__o211a_1 _6034_ (.A1(\core_0.execute.rf.reg_outputs[5][13] ),
    .A2(_2751_),
    .B1(_2758_),
    .C1(_2753_),
    .X(_0318_));
 sky130_fd_sc_hd__nand2_1 _6035_ (.A(_2713_),
    .B(_2742_),
    .Y(_2759_));
 sky130_fd_sc_hd__o211a_1 _6036_ (.A1(\core_0.execute.rf.reg_outputs[5][14] ),
    .A2(_2751_),
    .B1(_2759_),
    .C1(_2753_),
    .X(_0319_));
 sky130_fd_sc_hd__nand2_1 _6037_ (.A(_2716_),
    .B(_2742_),
    .Y(_2760_));
 sky130_fd_sc_hd__o211a_1 _6038_ (.A1(\core_0.execute.rf.reg_outputs[5][15] ),
    .A2(_2751_),
    .B1(_2760_),
    .C1(_2753_),
    .X(_0320_));
 sky130_fd_sc_hd__nand2_4 _6039_ (.A(\core_0.ew_reg_ie[4] ),
    .B(_2656_),
    .Y(_2761_));
 sky130_fd_sc_hd__and2_2 _6040_ (.A(\core_0.ew_reg_ie[4] ),
    .B(_2655_),
    .X(_2762_));
 sky130_fd_sc_hd__clkbuf_4 _6041_ (.A(_2762_),
    .X(_2763_));
 sky130_fd_sc_hd__or2_1 _6042_ (.A(\core_0.execute.rf.reg_outputs[4][0] ),
    .B(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__o211a_1 _6043_ (.A1(_2660_),
    .A2(_2761_),
    .B1(_2764_),
    .C1(_2753_),
    .X(_0321_));
 sky130_fd_sc_hd__or2_1 _6044_ (.A(\core_0.execute.rf.reg_outputs[4][1] ),
    .B(_2763_),
    .X(_2765_));
 sky130_fd_sc_hd__o211a_1 _6045_ (.A1(_2667_),
    .A2(_2761_),
    .B1(_2765_),
    .C1(_2753_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _6046_ (.A(\core_0.execute.rf.reg_outputs[4][2] ),
    .B(_2763_),
    .X(_2766_));
 sky130_fd_sc_hd__clkbuf_4 _6047_ (.A(_1314_),
    .X(_2767_));
 sky130_fd_sc_hd__o211a_1 _6048_ (.A1(_2671_),
    .A2(_2761_),
    .B1(_2766_),
    .C1(_2767_),
    .X(_0323_));
 sky130_fd_sc_hd__or2_1 _6049_ (.A(\core_0.execute.rf.reg_outputs[4][3] ),
    .B(_2763_),
    .X(_2768_));
 sky130_fd_sc_hd__o211a_1 _6050_ (.A1(_2675_),
    .A2(_2761_),
    .B1(_2768_),
    .C1(_2767_),
    .X(_0324_));
 sky130_fd_sc_hd__or2_1 _6051_ (.A(\core_0.execute.rf.reg_outputs[4][4] ),
    .B(_2762_),
    .X(_2769_));
 sky130_fd_sc_hd__o211a_1 _6052_ (.A1(_2679_),
    .A2(_2761_),
    .B1(_2769_),
    .C1(_2767_),
    .X(_0325_));
 sky130_fd_sc_hd__or2_1 _6053_ (.A(\core_0.execute.rf.reg_outputs[4][5] ),
    .B(_2762_),
    .X(_2770_));
 sky130_fd_sc_hd__o211a_1 _6054_ (.A1(_2683_),
    .A2(_2761_),
    .B1(_2770_),
    .C1(_2767_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_1 _6055_ (.A(\core_0.execute.rf.reg_outputs[4][6] ),
    .B(_2762_),
    .X(_2771_));
 sky130_fd_sc_hd__o211a_1 _6056_ (.A1(_2687_),
    .A2(_2761_),
    .B1(_2771_),
    .C1(_2767_),
    .X(_0327_));
 sky130_fd_sc_hd__or2_1 _6057_ (.A(\core_0.execute.rf.reg_outputs[4][7] ),
    .B(_2762_),
    .X(_2772_));
 sky130_fd_sc_hd__o211a_1 _6058_ (.A1(_2691_),
    .A2(_2761_),
    .B1(_2772_),
    .C1(_2767_),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_4 _6059_ (.A(_2762_),
    .X(_2773_));
 sky130_fd_sc_hd__nand2_1 _6060_ (.A(_2697_),
    .B(_2773_),
    .Y(_2774_));
 sky130_fd_sc_hd__o211a_1 _6061_ (.A1(\core_0.execute.rf.reg_outputs[4][8] ),
    .A2(_2773_),
    .B1(_2774_),
    .C1(_2767_),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_1 _6062_ (.A(_2699_),
    .B(_2773_),
    .Y(_2775_));
 sky130_fd_sc_hd__o211a_1 _6063_ (.A1(\core_0.execute.rf.reg_outputs[4][9] ),
    .A2(_2773_),
    .B1(_2775_),
    .C1(_2767_),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _6064_ (.A(_2701_),
    .B(_2763_),
    .Y(_2776_));
 sky130_fd_sc_hd__o211a_1 _6065_ (.A1(\core_0.execute.rf.reg_outputs[4][10] ),
    .A2(_2773_),
    .B1(_2776_),
    .C1(_2767_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_1 _6066_ (.A(_2705_),
    .B(_2763_),
    .Y(_2777_));
 sky130_fd_sc_hd__o211a_1 _6067_ (.A1(\core_0.execute.rf.reg_outputs[4][11] ),
    .A2(_2773_),
    .B1(_2777_),
    .C1(_2767_),
    .X(_0332_));
 sky130_fd_sc_hd__nand2_1 _6068_ (.A(_2707_),
    .B(_2763_),
    .Y(_2778_));
 sky130_fd_sc_hd__clkbuf_4 _6069_ (.A(_1314_),
    .X(_2779_));
 sky130_fd_sc_hd__o211a_1 _6070_ (.A1(\core_0.execute.rf.reg_outputs[4][12] ),
    .A2(_2773_),
    .B1(_2778_),
    .C1(_2779_),
    .X(_0333_));
 sky130_fd_sc_hd__nand2_1 _6071_ (.A(_2710_),
    .B(_2763_),
    .Y(_2780_));
 sky130_fd_sc_hd__o211a_1 _6072_ (.A1(\core_0.execute.rf.reg_outputs[4][13] ),
    .A2(_2773_),
    .B1(_2780_),
    .C1(_2779_),
    .X(_0334_));
 sky130_fd_sc_hd__nand2_1 _6073_ (.A(_2713_),
    .B(_2763_),
    .Y(_2781_));
 sky130_fd_sc_hd__o211a_1 _6074_ (.A1(\core_0.execute.rf.reg_outputs[4][14] ),
    .A2(_2773_),
    .B1(_2781_),
    .C1(_2779_),
    .X(_0335_));
 sky130_fd_sc_hd__nand2_1 _6075_ (.A(_2716_),
    .B(_2763_),
    .Y(_2782_));
 sky130_fd_sc_hd__o211a_1 _6076_ (.A1(\core_0.execute.rf.reg_outputs[4][15] ),
    .A2(_2773_),
    .B1(_2782_),
    .C1(_2779_),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_4 _6077_ (.A(\core_0.ew_reg_ie[3] ),
    .B(_2656_),
    .Y(_2783_));
 sky130_fd_sc_hd__and2_2 _6078_ (.A(\core_0.ew_reg_ie[3] ),
    .B(_2655_),
    .X(_2784_));
 sky130_fd_sc_hd__buf_2 _6079_ (.A(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__or2_1 _6080_ (.A(\core_0.execute.rf.reg_outputs[3][0] ),
    .B(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__o211a_1 _6081_ (.A1(_2660_),
    .A2(_2783_),
    .B1(_2786_),
    .C1(_2779_),
    .X(_0337_));
 sky130_fd_sc_hd__or2_1 _6082_ (.A(\core_0.execute.rf.reg_outputs[3][1] ),
    .B(_2785_),
    .X(_2787_));
 sky130_fd_sc_hd__o211a_1 _6083_ (.A1(_2667_),
    .A2(_2783_),
    .B1(_2787_),
    .C1(_2779_),
    .X(_0338_));
 sky130_fd_sc_hd__or2_1 _6084_ (.A(\core_0.execute.rf.reg_outputs[3][2] ),
    .B(_2785_),
    .X(_2788_));
 sky130_fd_sc_hd__o211a_1 _6085_ (.A1(_2671_),
    .A2(_2783_),
    .B1(_2788_),
    .C1(_2779_),
    .X(_0339_));
 sky130_fd_sc_hd__or2_1 _6086_ (.A(\core_0.execute.rf.reg_outputs[3][3] ),
    .B(_2785_),
    .X(_2789_));
 sky130_fd_sc_hd__o211a_1 _6087_ (.A1(_2675_),
    .A2(_2783_),
    .B1(_2789_),
    .C1(_2779_),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _6088_ (.A(\core_0.execute.rf.reg_outputs[3][4] ),
    .B(_2784_),
    .X(_2790_));
 sky130_fd_sc_hd__o211a_1 _6089_ (.A1(_2679_),
    .A2(_2783_),
    .B1(_2790_),
    .C1(_2779_),
    .X(_0341_));
 sky130_fd_sc_hd__or2_1 _6090_ (.A(\core_0.execute.rf.reg_outputs[3][5] ),
    .B(_2784_),
    .X(_2791_));
 sky130_fd_sc_hd__o211a_1 _6091_ (.A1(_2683_),
    .A2(_2783_),
    .B1(_2791_),
    .C1(_2779_),
    .X(_0342_));
 sky130_fd_sc_hd__or2_1 _6092_ (.A(\core_0.execute.rf.reg_outputs[3][6] ),
    .B(_2784_),
    .X(_2792_));
 sky130_fd_sc_hd__clkbuf_4 _6093_ (.A(_0996_),
    .X(_2793_));
 sky130_fd_sc_hd__o211a_1 _6094_ (.A1(_2687_),
    .A2(_2783_),
    .B1(_2792_),
    .C1(_2793_),
    .X(_0343_));
 sky130_fd_sc_hd__or2_1 _6095_ (.A(\core_0.execute.rf.reg_outputs[3][7] ),
    .B(_2784_),
    .X(_2794_));
 sky130_fd_sc_hd__o211a_1 _6096_ (.A1(_2691_),
    .A2(_2783_),
    .B1(_2794_),
    .C1(_2793_),
    .X(_0344_));
 sky130_fd_sc_hd__buf_2 _6097_ (.A(_2784_),
    .X(_2795_));
 sky130_fd_sc_hd__nand2_1 _6098_ (.A(_2697_),
    .B(_2795_),
    .Y(_2796_));
 sky130_fd_sc_hd__o211a_1 _6099_ (.A1(\core_0.execute.rf.reg_outputs[3][8] ),
    .A2(_2795_),
    .B1(_2796_),
    .C1(_2793_),
    .X(_0345_));
 sky130_fd_sc_hd__nand2_1 _6100_ (.A(_2699_),
    .B(_2795_),
    .Y(_2797_));
 sky130_fd_sc_hd__o211a_1 _6101_ (.A1(\core_0.execute.rf.reg_outputs[3][9] ),
    .A2(_2795_),
    .B1(_2797_),
    .C1(_2793_),
    .X(_0346_));
 sky130_fd_sc_hd__nand2_1 _6102_ (.A(_2701_),
    .B(_2785_),
    .Y(_2798_));
 sky130_fd_sc_hd__o211a_1 _6103_ (.A1(\core_0.execute.rf.reg_outputs[3][10] ),
    .A2(_2795_),
    .B1(_2798_),
    .C1(_2793_),
    .X(_0347_));
 sky130_fd_sc_hd__nand2_1 _6104_ (.A(_2705_),
    .B(_2785_),
    .Y(_2799_));
 sky130_fd_sc_hd__o211a_1 _6105_ (.A1(\core_0.execute.rf.reg_outputs[3][11] ),
    .A2(_2795_),
    .B1(_2799_),
    .C1(_2793_),
    .X(_0348_));
 sky130_fd_sc_hd__nand2_1 _6106_ (.A(_2707_),
    .B(_2785_),
    .Y(_2800_));
 sky130_fd_sc_hd__o211a_1 _6107_ (.A1(\core_0.execute.rf.reg_outputs[3][12] ),
    .A2(_2795_),
    .B1(_2800_),
    .C1(_2793_),
    .X(_0349_));
 sky130_fd_sc_hd__nand2_1 _6108_ (.A(_2710_),
    .B(_2785_),
    .Y(_2801_));
 sky130_fd_sc_hd__o211a_1 _6109_ (.A1(\core_0.execute.rf.reg_outputs[3][13] ),
    .A2(_2795_),
    .B1(_2801_),
    .C1(_2793_),
    .X(_0350_));
 sky130_fd_sc_hd__nand2_1 _6110_ (.A(_2713_),
    .B(_2785_),
    .Y(_2802_));
 sky130_fd_sc_hd__o211a_1 _6111_ (.A1(\core_0.execute.rf.reg_outputs[3][14] ),
    .A2(_2795_),
    .B1(_2802_),
    .C1(_2793_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_1 _6112_ (.A(_2716_),
    .B(_2785_),
    .Y(_2803_));
 sky130_fd_sc_hd__o211a_1 _6113_ (.A1(\core_0.execute.rf.reg_outputs[3][15] ),
    .A2(_2795_),
    .B1(_2803_),
    .C1(_2793_),
    .X(_0352_));
 sky130_fd_sc_hd__nand2_4 _6114_ (.A(\core_0.ew_reg_ie[2] ),
    .B(_2656_),
    .Y(_2804_));
 sky130_fd_sc_hd__and2_2 _6115_ (.A(\core_0.ew_reg_ie[2] ),
    .B(_2655_),
    .X(_2805_));
 sky130_fd_sc_hd__clkbuf_4 _6116_ (.A(_2805_),
    .X(_2806_));
 sky130_fd_sc_hd__or2_1 _6117_ (.A(\core_0.execute.rf.reg_outputs[2][0] ),
    .B(_2806_),
    .X(_2807_));
 sky130_fd_sc_hd__clkbuf_4 _6118_ (.A(_0996_),
    .X(_2808_));
 sky130_fd_sc_hd__o211a_1 _6119_ (.A1(_2660_),
    .A2(_2804_),
    .B1(_2807_),
    .C1(_2808_),
    .X(_0353_));
 sky130_fd_sc_hd__or2_1 _6120_ (.A(\core_0.execute.rf.reg_outputs[2][1] ),
    .B(_2806_),
    .X(_2809_));
 sky130_fd_sc_hd__o211a_1 _6121_ (.A1(_2667_),
    .A2(_2804_),
    .B1(_2809_),
    .C1(_2808_),
    .X(_0354_));
 sky130_fd_sc_hd__or2_1 _6122_ (.A(\core_0.execute.rf.reg_outputs[2][2] ),
    .B(_2806_),
    .X(_2810_));
 sky130_fd_sc_hd__o211a_1 _6123_ (.A1(_2671_),
    .A2(_2804_),
    .B1(_2810_),
    .C1(_2808_),
    .X(_0355_));
 sky130_fd_sc_hd__or2_1 _6124_ (.A(\core_0.execute.rf.reg_outputs[2][3] ),
    .B(_2806_),
    .X(_2811_));
 sky130_fd_sc_hd__o211a_1 _6125_ (.A1(_2675_),
    .A2(_2804_),
    .B1(_2811_),
    .C1(_2808_),
    .X(_0356_));
 sky130_fd_sc_hd__or2_1 _6126_ (.A(\core_0.execute.rf.reg_outputs[2][4] ),
    .B(_2805_),
    .X(_2812_));
 sky130_fd_sc_hd__o211a_1 _6127_ (.A1(_2679_),
    .A2(_2804_),
    .B1(_2812_),
    .C1(_2808_),
    .X(_0357_));
 sky130_fd_sc_hd__or2_1 _6128_ (.A(\core_0.execute.rf.reg_outputs[2][5] ),
    .B(_2805_),
    .X(_2813_));
 sky130_fd_sc_hd__o211a_1 _6129_ (.A1(_2683_),
    .A2(_2804_),
    .B1(_2813_),
    .C1(_2808_),
    .X(_0358_));
 sky130_fd_sc_hd__or2_1 _6130_ (.A(\core_0.execute.rf.reg_outputs[2][6] ),
    .B(_2805_),
    .X(_2814_));
 sky130_fd_sc_hd__o211a_1 _6131_ (.A1(_2687_),
    .A2(_2804_),
    .B1(_2814_),
    .C1(_2808_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _6132_ (.A(\core_0.execute.rf.reg_outputs[2][7] ),
    .B(_2805_),
    .X(_2815_));
 sky130_fd_sc_hd__o211a_1 _6133_ (.A1(_2691_),
    .A2(_2804_),
    .B1(_2815_),
    .C1(_2808_),
    .X(_0360_));
 sky130_fd_sc_hd__buf_2 _6134_ (.A(_2805_),
    .X(_2816_));
 sky130_fd_sc_hd__nand2_1 _6135_ (.A(_2697_),
    .B(_2816_),
    .Y(_2817_));
 sky130_fd_sc_hd__o211a_1 _6136_ (.A1(\core_0.execute.rf.reg_outputs[2][8] ),
    .A2(_2816_),
    .B1(_2817_),
    .C1(_2808_),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_1 _6137_ (.A(_2699_),
    .B(_2816_),
    .Y(_2818_));
 sky130_fd_sc_hd__o211a_1 _6138_ (.A1(\core_0.execute.rf.reg_outputs[2][9] ),
    .A2(_2816_),
    .B1(_2818_),
    .C1(_2808_),
    .X(_0362_));
 sky130_fd_sc_hd__nand2_1 _6139_ (.A(_2701_),
    .B(_2806_),
    .Y(_2819_));
 sky130_fd_sc_hd__clkbuf_4 _6140_ (.A(_0996_),
    .X(_2820_));
 sky130_fd_sc_hd__o211a_1 _6141_ (.A1(\core_0.execute.rf.reg_outputs[2][10] ),
    .A2(_2816_),
    .B1(_2819_),
    .C1(_2820_),
    .X(_0363_));
 sky130_fd_sc_hd__nand2_1 _6142_ (.A(_2705_),
    .B(_2806_),
    .Y(_2821_));
 sky130_fd_sc_hd__o211a_1 _6143_ (.A1(\core_0.execute.rf.reg_outputs[2][11] ),
    .A2(_2816_),
    .B1(_2821_),
    .C1(_2820_),
    .X(_0364_));
 sky130_fd_sc_hd__nand2_1 _6144_ (.A(_2707_),
    .B(_2806_),
    .Y(_2822_));
 sky130_fd_sc_hd__o211a_1 _6145_ (.A1(\core_0.execute.rf.reg_outputs[2][12] ),
    .A2(_2816_),
    .B1(_2822_),
    .C1(_2820_),
    .X(_0365_));
 sky130_fd_sc_hd__nand2_1 _6146_ (.A(_2710_),
    .B(_2806_),
    .Y(_2823_));
 sky130_fd_sc_hd__o211a_1 _6147_ (.A1(\core_0.execute.rf.reg_outputs[2][13] ),
    .A2(_2816_),
    .B1(_2823_),
    .C1(_2820_),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_1 _6148_ (.A(_2713_),
    .B(_2806_),
    .Y(_2824_));
 sky130_fd_sc_hd__o211a_1 _6149_ (.A1(\core_0.execute.rf.reg_outputs[2][14] ),
    .A2(_2816_),
    .B1(_2824_),
    .C1(_2820_),
    .X(_0367_));
 sky130_fd_sc_hd__nand2_1 _6150_ (.A(_2716_),
    .B(_2806_),
    .Y(_2825_));
 sky130_fd_sc_hd__o211a_1 _6151_ (.A1(\core_0.execute.rf.reg_outputs[2][15] ),
    .A2(_2816_),
    .B1(_2825_),
    .C1(_2820_),
    .X(_0368_));
 sky130_fd_sc_hd__nand2_4 _6152_ (.A(\core_0.ew_reg_ie[1] ),
    .B(_2656_),
    .Y(_2826_));
 sky130_fd_sc_hd__and2_1 _6153_ (.A(\core_0.ew_reg_ie[1] ),
    .B(_2655_),
    .X(_2827_));
 sky130_fd_sc_hd__clkbuf_4 _6154_ (.A(_2827_),
    .X(_2828_));
 sky130_fd_sc_hd__or2_1 _6155_ (.A(\core_0.execute.rf.reg_outputs[1][0] ),
    .B(_2828_),
    .X(_2829_));
 sky130_fd_sc_hd__o211a_1 _6156_ (.A1(_2660_),
    .A2(_2826_),
    .B1(_2829_),
    .C1(_2820_),
    .X(_0369_));
 sky130_fd_sc_hd__or2_1 _6157_ (.A(\core_0.execute.rf.reg_outputs[1][1] ),
    .B(_2828_),
    .X(_2830_));
 sky130_fd_sc_hd__o211a_1 _6158_ (.A1(_2667_),
    .A2(_2826_),
    .B1(_2830_),
    .C1(_2820_),
    .X(_0370_));
 sky130_fd_sc_hd__or2_1 _6159_ (.A(\core_0.execute.rf.reg_outputs[1][2] ),
    .B(_2828_),
    .X(_2831_));
 sky130_fd_sc_hd__o211a_1 _6160_ (.A1(_2671_),
    .A2(_2826_),
    .B1(_2831_),
    .C1(_2820_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _6161_ (.A(\core_0.execute.rf.reg_outputs[1][3] ),
    .B(_2828_),
    .X(_2832_));
 sky130_fd_sc_hd__o211a_1 _6162_ (.A1(_2675_),
    .A2(_2826_),
    .B1(_2832_),
    .C1(_2820_),
    .X(_0372_));
 sky130_fd_sc_hd__or2_1 _6163_ (.A(\core_0.execute.rf.reg_outputs[1][4] ),
    .B(_2827_),
    .X(_2833_));
 sky130_fd_sc_hd__buf_4 _6164_ (.A(_0996_),
    .X(_2834_));
 sky130_fd_sc_hd__o211a_1 _6165_ (.A1(_2679_),
    .A2(_2826_),
    .B1(_2833_),
    .C1(_2834_),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _6166_ (.A(\core_0.execute.rf.reg_outputs[1][5] ),
    .B(_2827_),
    .X(_2835_));
 sky130_fd_sc_hd__o211a_1 _6167_ (.A1(_2683_),
    .A2(_2826_),
    .B1(_2835_),
    .C1(_2834_),
    .X(_0374_));
 sky130_fd_sc_hd__or2_1 _6168_ (.A(\core_0.execute.rf.reg_outputs[1][6] ),
    .B(_2827_),
    .X(_2836_));
 sky130_fd_sc_hd__o211a_1 _6169_ (.A1(_2687_),
    .A2(_2826_),
    .B1(_2836_),
    .C1(_2834_),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _6170_ (.A(\core_0.execute.rf.reg_outputs[1][7] ),
    .B(_2827_),
    .X(_2837_));
 sky130_fd_sc_hd__o211a_1 _6171_ (.A1(_2691_),
    .A2(_2826_),
    .B1(_2837_),
    .C1(_2834_),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_4 _6172_ (.A(_2827_),
    .X(_2838_));
 sky130_fd_sc_hd__nand2_1 _6173_ (.A(_2697_),
    .B(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__o211a_1 _6174_ (.A1(\core_0.execute.rf.reg_outputs[1][8] ),
    .A2(_2838_),
    .B1(_2839_),
    .C1(_2834_),
    .X(_0377_));
 sky130_fd_sc_hd__nand2_1 _6175_ (.A(_2699_),
    .B(_2838_),
    .Y(_2840_));
 sky130_fd_sc_hd__o211a_1 _6176_ (.A1(\core_0.execute.rf.reg_outputs[1][9] ),
    .A2(_2838_),
    .B1(_2840_),
    .C1(_2834_),
    .X(_0378_));
 sky130_fd_sc_hd__nand2_1 _6177_ (.A(_2701_),
    .B(_2828_),
    .Y(_2841_));
 sky130_fd_sc_hd__o211a_1 _6178_ (.A1(\core_0.execute.rf.reg_outputs[1][10] ),
    .A2(_2838_),
    .B1(_2841_),
    .C1(_2834_),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_1 _6179_ (.A(_2705_),
    .B(_2828_),
    .Y(_2842_));
 sky130_fd_sc_hd__o211a_1 _6180_ (.A1(\core_0.execute.rf.reg_outputs[1][11] ),
    .A2(_2838_),
    .B1(_2842_),
    .C1(_2834_),
    .X(_0380_));
 sky130_fd_sc_hd__nand2_1 _6181_ (.A(_2707_),
    .B(_2828_),
    .Y(_2843_));
 sky130_fd_sc_hd__o211a_1 _6182_ (.A1(\core_0.execute.rf.reg_outputs[1][12] ),
    .A2(_2838_),
    .B1(_2843_),
    .C1(_2834_),
    .X(_0381_));
 sky130_fd_sc_hd__nand2_1 _6183_ (.A(_2710_),
    .B(_2828_),
    .Y(_2844_));
 sky130_fd_sc_hd__o211a_1 _6184_ (.A1(\core_0.execute.rf.reg_outputs[1][13] ),
    .A2(_2838_),
    .B1(_2844_),
    .C1(_2834_),
    .X(_0382_));
 sky130_fd_sc_hd__nand2_1 _6185_ (.A(_2713_),
    .B(_2828_),
    .Y(_2845_));
 sky130_fd_sc_hd__buf_2 _6186_ (.A(_0996_),
    .X(_2846_));
 sky130_fd_sc_hd__o211a_1 _6187_ (.A1(\core_0.execute.rf.reg_outputs[1][14] ),
    .A2(_2838_),
    .B1(_2845_),
    .C1(_2846_),
    .X(_0383_));
 sky130_fd_sc_hd__nand2_1 _6188_ (.A(_2716_),
    .B(_2828_),
    .Y(_2847_));
 sky130_fd_sc_hd__o211a_1 _6189_ (.A1(\core_0.execute.rf.reg_outputs[1][15] ),
    .A2(_2838_),
    .B1(_2847_),
    .C1(_2846_),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_2 _6190_ (.A(\core_0.ew_reg_ie[0] ),
    .B(_2656_),
    .Y(_2848_));
 sky130_fd_sc_hd__and2_1 _6191_ (.A(\core_0.ew_reg_ie[0] ),
    .B(_2655_),
    .X(_2849_));
 sky130_fd_sc_hd__buf_2 _6192_ (.A(_2849_),
    .X(_2850_));
 sky130_fd_sc_hd__or2_1 _6193_ (.A(net88),
    .B(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__o211a_1 _6194_ (.A1(_2660_),
    .A2(_2848_),
    .B1(_2851_),
    .C1(_2846_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _6195_ (.A(net95),
    .B(_2850_),
    .X(_2852_));
 sky130_fd_sc_hd__o211a_1 _6196_ (.A1(_2667_),
    .A2(_2848_),
    .B1(_2852_),
    .C1(_2846_),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _6197_ (.A(net96),
    .B(_2850_),
    .X(_2853_));
 sky130_fd_sc_hd__o211a_1 _6198_ (.A1(_2671_),
    .A2(_2848_),
    .B1(_2853_),
    .C1(_2846_),
    .X(_0387_));
 sky130_fd_sc_hd__or2_1 _6199_ (.A(net97),
    .B(_2850_),
    .X(_2854_));
 sky130_fd_sc_hd__o211a_1 _6200_ (.A1(_2675_),
    .A2(_2848_),
    .B1(_2854_),
    .C1(_2846_),
    .X(_0388_));
 sky130_fd_sc_hd__or2_1 _6201_ (.A(net98),
    .B(_2849_),
    .X(_2855_));
 sky130_fd_sc_hd__o211a_1 _6202_ (.A1(_2679_),
    .A2(_2848_),
    .B1(_2855_),
    .C1(_2846_),
    .X(_0389_));
 sky130_fd_sc_hd__or2_1 _6203_ (.A(net99),
    .B(_2849_),
    .X(_2856_));
 sky130_fd_sc_hd__o211a_1 _6204_ (.A1(_2683_),
    .A2(_2848_),
    .B1(_2856_),
    .C1(_2846_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_1 _6205_ (.A(net100),
    .B(_2849_),
    .X(_2857_));
 sky130_fd_sc_hd__o211a_1 _6206_ (.A1(_2687_),
    .A2(_2848_),
    .B1(_2857_),
    .C1(_2846_),
    .X(_0391_));
 sky130_fd_sc_hd__or2_1 _6207_ (.A(net101),
    .B(_2849_),
    .X(_2858_));
 sky130_fd_sc_hd__o211a_1 _6208_ (.A1(_2691_),
    .A2(_2848_),
    .B1(_2858_),
    .C1(_2846_),
    .X(_0392_));
 sky130_fd_sc_hd__buf_2 _6209_ (.A(_2849_),
    .X(_2859_));
 sky130_fd_sc_hd__nand2_1 _6210_ (.A(_2697_),
    .B(_2859_),
    .Y(_2860_));
 sky130_fd_sc_hd__buf_6 _6211_ (.A(_0996_),
    .X(_2861_));
 sky130_fd_sc_hd__o211a_1 _6212_ (.A1(net102),
    .A2(_2859_),
    .B1(_2860_),
    .C1(_2861_),
    .X(_0393_));
 sky130_fd_sc_hd__nand2_1 _6213_ (.A(_2699_),
    .B(_2859_),
    .Y(_2862_));
 sky130_fd_sc_hd__o211a_1 _6214_ (.A1(net103),
    .A2(_2859_),
    .B1(_2862_),
    .C1(_2861_),
    .X(_0394_));
 sky130_fd_sc_hd__nand2_1 _6215_ (.A(_2701_),
    .B(_2850_),
    .Y(_2863_));
 sky130_fd_sc_hd__o211a_1 _6216_ (.A1(net89),
    .A2(_2859_),
    .B1(_2863_),
    .C1(_2861_),
    .X(_0395_));
 sky130_fd_sc_hd__nand2_1 _6217_ (.A(_2705_),
    .B(_2850_),
    .Y(_2864_));
 sky130_fd_sc_hd__o211a_1 _6218_ (.A1(net90),
    .A2(_2859_),
    .B1(_2864_),
    .C1(_2861_),
    .X(_0396_));
 sky130_fd_sc_hd__nand2_1 _6219_ (.A(_2707_),
    .B(_2850_),
    .Y(_2865_));
 sky130_fd_sc_hd__o211a_1 _6220_ (.A1(net91),
    .A2(_2859_),
    .B1(_2865_),
    .C1(_2861_),
    .X(_0397_));
 sky130_fd_sc_hd__nand2_1 _6221_ (.A(_2710_),
    .B(_2850_),
    .Y(_2866_));
 sky130_fd_sc_hd__o211a_1 _6222_ (.A1(net92),
    .A2(_2859_),
    .B1(_2866_),
    .C1(_2861_),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_1 _6223_ (.A(_2713_),
    .B(_2850_),
    .Y(_2867_));
 sky130_fd_sc_hd__o211a_1 _6224_ (.A1(net93),
    .A2(_2859_),
    .B1(_2867_),
    .C1(_2861_),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_1 _6225_ (.A(_2716_),
    .B(_2850_),
    .Y(_2868_));
 sky130_fd_sc_hd__o211a_1 _6226_ (.A1(net94),
    .A2(_2859_),
    .B1(_2868_),
    .C1(_2861_),
    .X(_0400_));
 sky130_fd_sc_hd__nor2_1 _6227_ (.A(_0907_),
    .B(_0674_),
    .Y(_2869_));
 sky130_fd_sc_hd__buf_4 _6228_ (.A(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__a21oi_1 _6229_ (.A1(_1154_),
    .A2(_1027_),
    .B1(\core_0.execute.irq_en ),
    .Y(_2871_));
 sky130_fd_sc_hd__nand2_1 _6230_ (.A(_1163_),
    .B(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__o211a_1 _6231_ (.A1(net202),
    .A2(_1169_),
    .B1(_2870_),
    .C1(_2872_),
    .X(_0401_));
 sky130_fd_sc_hd__and2_1 _6232_ (.A(\core_0.decode.o_submit ),
    .B(_0955_),
    .X(_2873_));
 sky130_fd_sc_hd__buf_2 _6233_ (.A(_2873_),
    .X(_2874_));
 sky130_fd_sc_hd__clkbuf_4 _6234_ (.A(_2874_),
    .X(_2875_));
 sky130_fd_sc_hd__a211o_1 _6235_ (.A1(_1560_),
    .A2(_0742_),
    .B1(_2875_),
    .C1(_1795_),
    .X(_2876_));
 sky130_fd_sc_hd__o21a_1 _6236_ (.A1(_1205_),
    .A2(_1212_),
    .B1(_2876_),
    .X(_0402_));
 sky130_fd_sc_hd__nand2_1 _6237_ (.A(_1560_),
    .B(_1207_),
    .Y(_2877_));
 sky130_fd_sc_hd__nor2_1 _6238_ (.A(_1344_),
    .B(_2877_),
    .Y(_2878_));
 sky130_fd_sc_hd__a221o_1 _6239_ (.A1(_1437_),
    .A2(_1342_),
    .B1(_1350_),
    .B2(_1602_),
    .C1(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__a211oi_2 _6240_ (.A1(_1797_),
    .A2(_1392_),
    .B1(_2879_),
    .C1(_1436_),
    .Y(_2880_));
 sky130_fd_sc_hd__nand2_1 _6241_ (.A(_1334_),
    .B(_1602_),
    .Y(_2881_));
 sky130_fd_sc_hd__o221a_1 _6242_ (.A1(_1603_),
    .A2(_1400_),
    .B1(_2877_),
    .B2(_1331_),
    .C1(_2881_),
    .X(_2882_));
 sky130_fd_sc_hd__o211a_1 _6243_ (.A1(_1208_),
    .A2(_1839_),
    .B1(_2882_),
    .C1(_1436_),
    .X(_2883_));
 sky130_fd_sc_hd__nand2_1 _6244_ (.A(_1362_),
    .B(_1602_),
    .Y(_2884_));
 sky130_fd_sc_hd__o221a_1 _6245_ (.A1(_1603_),
    .A2(_1701_),
    .B1(_2877_),
    .B2(_1357_),
    .C1(_2884_),
    .X(_2885_));
 sky130_fd_sc_hd__o211a_1 _6246_ (.A1(_1208_),
    .A2(_1902_),
    .B1(_2885_),
    .C1(_1435_),
    .X(_2886_));
 sky130_fd_sc_hd__nand2_1 _6247_ (.A(_1739_),
    .B(_1602_),
    .Y(_2887_));
 sky130_fd_sc_hd__o221a_1 _6248_ (.A1(_1603_),
    .A2(_2002_),
    .B1(_2877_),
    .B2(_1749_),
    .C1(_2887_),
    .X(_2888_));
 sky130_fd_sc_hd__o211a_1 _6249_ (.A1(_1208_),
    .A2(_1751_),
    .B1(_2888_),
    .C1(_1204_),
    .X(_2889_));
 sky130_fd_sc_hd__o311a_1 _6250_ (.A1(_1202_),
    .A2(_2886_),
    .A3(_2889_),
    .B1(\core_0.execute.alu_mul_div.comp ),
    .C1(_0955_),
    .X(_2890_));
 sky130_fd_sc_hd__o31ai_4 _6251_ (.A1(_1803_),
    .A2(_2880_),
    .A3(_2883_),
    .B1(_2890_),
    .Y(_2891_));
 sky130_fd_sc_hd__nor2_4 _6252_ (.A(\core_0.decode.o_submit ),
    .B(_2891_),
    .Y(_2892_));
 sky130_fd_sc_hd__and3_1 _6253_ (.A(_1802_),
    .B(_1203_),
    .C(_1797_),
    .X(_2893_));
 sky130_fd_sc_hd__and3_1 _6254_ (.A(\core_0.execute.alu_mul_div.mul_res[0] ),
    .B(_1644_),
    .C(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__a21oi_1 _6255_ (.A1(_1644_),
    .A2(_2893_),
    .B1(\core_0.execute.alu_mul_div.mul_res[0] ),
    .Y(_2895_));
 sky130_fd_sc_hd__nor2_1 _6256_ (.A(_2894_),
    .B(_2895_),
    .Y(_2896_));
 sky130_fd_sc_hd__and2_2 _6257_ (.A(_0743_),
    .B(_2891_),
    .X(_2897_));
 sky130_fd_sc_hd__clkbuf_4 _6258_ (.A(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__a22o_1 _6259_ (.A1(_2892_),
    .A2(_2896_),
    .B1(_2898_),
    .B2(\core_0.execute.alu_mul_div.mul_res[0] ),
    .X(_2899_));
 sky130_fd_sc_hd__a21o_1 _6260_ (.A1(_2875_),
    .A2(_1767_),
    .B1(_2899_),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_4 _6261_ (.A(_2002_),
    .X(_2900_));
 sky130_fd_sc_hd__and4_4 _6262_ (.A(_1559_),
    .B(_1617_),
    .C(_1621_),
    .D(_1622_),
    .X(_2901_));
 sky130_fd_sc_hd__a2111oi_4 _6263_ (.A1(_1205_),
    .A2(_1766_),
    .B1(_2901_),
    .C1(\core_0.execute.alu_mul_div.cbit[1] ),
    .D1(\core_0.execute.alu_mul_div.cbit[2] ),
    .Y(_2902_));
 sky130_fd_sc_hd__and3_1 _6264_ (.A(_1802_),
    .B(\core_0.execute.alu_mul_div.mul_res[1] ),
    .C(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__a21o_1 _6265_ (.A1(_1802_),
    .A2(_2902_),
    .B1(\core_0.execute.alu_mul_div.mul_res[1] ),
    .X(_2904_));
 sky130_fd_sc_hd__or2b_1 _6266_ (.A(_2903_),
    .B_N(_2904_),
    .X(_2905_));
 sky130_fd_sc_hd__xnor2_1 _6267_ (.A(_2894_),
    .B(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__a22o_1 _6268_ (.A1(\core_0.execute.alu_mul_div.mul_res[1] ),
    .A2(_2898_),
    .B1(_2906_),
    .B2(_2892_),
    .X(_2907_));
 sky130_fd_sc_hd__a31o_1 _6269_ (.A1(_2875_),
    .A2(_2900_),
    .A3(_1732_),
    .B1(_2907_),
    .X(_0404_));
 sky130_fd_sc_hd__and4_1 _6270_ (.A(_1802_),
    .B(_1203_),
    .C(\core_0.execute.alu_mul_div.mul_res[2] ),
    .D(_1646_),
    .X(_2908_));
 sky130_fd_sc_hd__a31o_1 _6271_ (.A1(_1802_),
    .A2(_1203_),
    .A3(_1646_),
    .B1(\core_0.execute.alu_mul_div.mul_res[2] ),
    .X(_2909_));
 sky130_fd_sc_hd__or2b_1 _6272_ (.A(_2908_),
    .B_N(_2909_),
    .X(_2910_));
 sky130_fd_sc_hd__a21o_1 _6273_ (.A1(_2894_),
    .A2(_2904_),
    .B1(_2903_),
    .X(_2911_));
 sky130_fd_sc_hd__xnor2_1 _6274_ (.A(_2910_),
    .B(_2911_),
    .Y(_2912_));
 sky130_fd_sc_hd__a22o_1 _6275_ (.A1(_2875_),
    .A2(_2128_),
    .B1(_2898_),
    .B2(\core_0.execute.alu_mul_div.mul_res[2] ),
    .X(_2913_));
 sky130_fd_sc_hd__a21o_1 _6276_ (.A1(_2892_),
    .A2(_2912_),
    .B1(_2913_),
    .X(_0405_));
 sky130_fd_sc_hd__mux4_2 _6277_ (.A0(_1633_),
    .A1(_1670_),
    .A2(_1766_),
    .A3(_1624_),
    .S0(_1559_),
    .S1(\core_0.execute.alu_mul_div.cbit[1] ),
    .X(_2914_));
 sky130_fd_sc_hd__or3_1 _6278_ (.A(\core_0.execute.alu_mul_div.cbit[3] ),
    .B(\core_0.execute.alu_mul_div.cbit[2] ),
    .C(_2914_),
    .X(_2915_));
 sky130_fd_sc_hd__xor2_1 _6279_ (.A(\core_0.execute.alu_mul_div.mul_res[3] ),
    .B(_2915_),
    .X(_2916_));
 sky130_fd_sc_hd__a21oi_1 _6280_ (.A1(_2909_),
    .A2(_2911_),
    .B1(_2908_),
    .Y(_2917_));
 sky130_fd_sc_hd__or2_1 _6281_ (.A(_2916_),
    .B(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__a21oi_1 _6282_ (.A1(_2916_),
    .A2(_2917_),
    .B1(_2874_),
    .Y(_2919_));
 sky130_fd_sc_hd__a32o_1 _6283_ (.A1(_2874_),
    .A2(_2900_),
    .A3(_2231_),
    .B1(_2918_),
    .B2(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__mux2_1 _6284_ (.A0(_2920_),
    .A1(\core_0.execute.alu_mul_div.mul_res[3] ),
    .S(_2898_),
    .X(_2921_));
 sky130_fd_sc_hd__clkbuf_1 _6285_ (.A(_2921_),
    .X(_0406_));
 sky130_fd_sc_hd__nand2_1 _6286_ (.A(_1797_),
    .B(_1644_),
    .Y(_2922_));
 sky130_fd_sc_hd__mux2_1 _6287_ (.A0(_1678_),
    .A1(_1634_),
    .S(_1206_),
    .X(_2923_));
 sky130_fd_sc_hd__mux2_1 _6288_ (.A0(_2922_),
    .A1(_2923_),
    .S(_1203_),
    .X(_2924_));
 sky130_fd_sc_hd__nor3b_1 _6289_ (.A(_1201_),
    .B(_2924_),
    .C_N(\core_0.execute.alu_mul_div.mul_res[4] ),
    .Y(_2925_));
 sky130_fd_sc_hd__o21ba_1 _6290_ (.A1(_1201_),
    .A2(_2924_),
    .B1_N(\core_0.execute.alu_mul_div.mul_res[4] ),
    .X(_2926_));
 sky130_fd_sc_hd__or2_1 _6291_ (.A(_2925_),
    .B(_2926_),
    .X(_2927_));
 sky130_fd_sc_hd__or2_1 _6292_ (.A(\core_0.execute.alu_mul_div.cbit[2] ),
    .B(_2914_),
    .X(_2928_));
 sky130_fd_sc_hd__or3b_1 _6293_ (.A(_2928_),
    .B(_1201_),
    .C_N(\core_0.execute.alu_mul_div.mul_res[3] ),
    .X(_2929_));
 sky130_fd_sc_hd__o21a_1 _6294_ (.A1(_2916_),
    .A2(_2917_),
    .B1(_2929_),
    .X(_2930_));
 sky130_fd_sc_hd__and2_1 _6295_ (.A(_2927_),
    .B(_2930_),
    .X(_2931_));
 sky130_fd_sc_hd__o21ai_1 _6296_ (.A1(_2927_),
    .A2(_2930_),
    .B1(_0743_),
    .Y(_2932_));
 sky130_fd_sc_hd__o22ai_1 _6297_ (.A1(_0743_),
    .A2(_2126_),
    .B1(_2931_),
    .B2(_2932_),
    .Y(_2933_));
 sky130_fd_sc_hd__mux2_1 _6298_ (.A0(_2933_),
    .A1(\core_0.execute.alu_mul_div.mul_res[4] ),
    .S(_2897_),
    .X(_2934_));
 sky130_fd_sc_hd__clkbuf_1 _6299_ (.A(_2934_),
    .X(_0407_));
 sky130_fd_sc_hd__nor2_1 _6300_ (.A(_1560_),
    .B(_1644_),
    .Y(_2935_));
 sky130_fd_sc_hd__mux4_1 _6301_ (.A0(_1743_),
    .A1(_1670_),
    .A2(_1677_),
    .A3(_1633_),
    .S0(\core_0.execute.alu_mul_div.cbit[1] ),
    .S1(_1205_),
    .X(_2936_));
 sky130_fd_sc_hd__or2_1 _6302_ (.A(\core_0.execute.alu_mul_div.cbit[2] ),
    .B(_2936_),
    .X(_2937_));
 sky130_fd_sc_hd__o41a_1 _6303_ (.A1(_1203_),
    .A2(_1206_),
    .A3(_2901_),
    .A4(_2935_),
    .B1(_2937_),
    .X(_2938_));
 sky130_fd_sc_hd__or3b_1 _6304_ (.A(_2938_),
    .B(_1201_),
    .C_N(\core_0.execute.alu_mul_div.mul_res[5] ),
    .X(_2939_));
 sky130_fd_sc_hd__o21bai_1 _6305_ (.A1(_1201_),
    .A2(_2938_),
    .B1_N(\core_0.execute.alu_mul_div.mul_res[5] ),
    .Y(_2940_));
 sky130_fd_sc_hd__nand2_1 _6306_ (.A(_2939_),
    .B(_2940_),
    .Y(_2941_));
 sky130_fd_sc_hd__o21bai_1 _6307_ (.A1(_2926_),
    .A2(_2930_),
    .B1_N(_2925_),
    .Y(_2942_));
 sky130_fd_sc_hd__xnor2_1 _6308_ (.A(_2941_),
    .B(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__and3_1 _6309_ (.A(_2875_),
    .B(_2900_),
    .C(_1661_),
    .X(_2944_));
 sky130_fd_sc_hd__a221o_1 _6310_ (.A1(\core_0.execute.alu_mul_div.mul_res[5] ),
    .A2(_2898_),
    .B1(_2943_),
    .B2(_2892_),
    .C1(_2944_),
    .X(_0408_));
 sky130_fd_sc_hd__or3b_1 _6311_ (.A(_1680_),
    .B(_1201_),
    .C_N(\core_0.execute.alu_mul_div.mul_res[6] ),
    .X(_2945_));
 sky130_fd_sc_hd__a21o_1 _6312_ (.A1(_1802_),
    .A2(_1681_),
    .B1(\core_0.execute.alu_mul_div.mul_res[6] ),
    .X(_2946_));
 sky130_fd_sc_hd__nand2_1 _6313_ (.A(_2945_),
    .B(_2946_),
    .Y(_2947_));
 sky130_fd_sc_hd__a21bo_1 _6314_ (.A1(_2940_),
    .A2(_2942_),
    .B1_N(_2939_),
    .X(_2948_));
 sky130_fd_sc_hd__xnor2_1 _6315_ (.A(_2947_),
    .B(_2948_),
    .Y(_2949_));
 sky130_fd_sc_hd__and3_1 _6316_ (.A(_2874_),
    .B(_2002_),
    .C(_1654_),
    .X(_2950_));
 sky130_fd_sc_hd__a21o_1 _6317_ (.A1(_0743_),
    .A2(_2949_),
    .B1(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__inv_2 _6318_ (.A(_2897_),
    .Y(_2952_));
 sky130_fd_sc_hd__mux2_1 _6319_ (.A0(\core_0.execute.alu_mul_div.mul_res[6] ),
    .A1(_2951_),
    .S(_2952_),
    .X(_2953_));
 sky130_fd_sc_hd__clkbuf_1 _6320_ (.A(_2953_),
    .X(_0409_));
 sky130_fd_sc_hd__mux4_2 _6321_ (.A0(_1745_),
    .A1(_1746_),
    .A2(_1743_),
    .A3(_1677_),
    .S0(_1205_),
    .S1(_1206_),
    .X(_2954_));
 sky130_fd_sc_hd__mux2_1 _6322_ (.A0(_2914_),
    .A1(_2954_),
    .S(_1204_),
    .X(_2955_));
 sky130_fd_sc_hd__nor2_1 _6323_ (.A(_1201_),
    .B(_2955_),
    .Y(_2956_));
 sky130_fd_sc_hd__and2_1 _6324_ (.A(\core_0.execute.alu_mul_div.mul_res[7] ),
    .B(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__nor2_1 _6325_ (.A(\core_0.execute.alu_mul_div.mul_res[7] ),
    .B(_2956_),
    .Y(_2958_));
 sky130_fd_sc_hd__or2_1 _6326_ (.A(_2957_),
    .B(_2958_),
    .X(_2959_));
 sky130_fd_sc_hd__a21boi_1 _6327_ (.A1(_2946_),
    .A2(_2948_),
    .B1_N(_2945_),
    .Y(_2960_));
 sky130_fd_sc_hd__nor2_1 _6328_ (.A(_2959_),
    .B(_2960_),
    .Y(_2961_));
 sky130_fd_sc_hd__inv_2 _6329_ (.A(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__nand2_1 _6330_ (.A(_2959_),
    .B(_2960_),
    .Y(_2963_));
 sky130_fd_sc_hd__a32o_1 _6331_ (.A1(_2875_),
    .A2(_2900_),
    .A3(_1571_),
    .B1(_2898_),
    .B2(\core_0.execute.alu_mul_div.mul_res[7] ),
    .X(_2964_));
 sky130_fd_sc_hd__a31o_1 _6332_ (.A1(_2892_),
    .A2(_2962_),
    .A3(_2963_),
    .B1(_2964_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _6333_ (.A0(_1580_),
    .A1(_1662_),
    .S(_1206_),
    .X(_2965_));
 sky130_fd_sc_hd__nor2_1 _6334_ (.A(\core_0.execute.alu_mul_div.cbit[2] ),
    .B(_2965_),
    .Y(_2966_));
 sky130_fd_sc_hd__a21o_1 _6335_ (.A1(\core_0.execute.alu_mul_div.cbit[2] ),
    .A2(_2923_),
    .B1(_1201_),
    .X(_2967_));
 sky130_fd_sc_hd__o32a_1 _6336_ (.A1(_1802_),
    .A2(_1435_),
    .A3(_2922_),
    .B1(_2966_),
    .B2(_2967_),
    .X(_2968_));
 sky130_fd_sc_hd__and2b_1 _6337_ (.A_N(_2968_),
    .B(\core_0.execute.alu_mul_div.mul_res[8] ),
    .X(_2969_));
 sky130_fd_sc_hd__and2b_1 _6338_ (.A_N(\core_0.execute.alu_mul_div.mul_res[8] ),
    .B(_2968_),
    .X(_2970_));
 sky130_fd_sc_hd__nor2_1 _6339_ (.A(_2969_),
    .B(_2970_),
    .Y(_2971_));
 sky130_fd_sc_hd__o21bai_1 _6340_ (.A1(_2959_),
    .A2(_2960_),
    .B1_N(_2957_),
    .Y(_2972_));
 sky130_fd_sc_hd__nand2_1 _6341_ (.A(_2971_),
    .B(_2972_),
    .Y(_2973_));
 sky130_fd_sc_hd__or2_1 _6342_ (.A(_2971_),
    .B(_2972_),
    .X(_2974_));
 sky130_fd_sc_hd__a31o_1 _6343_ (.A1(_2874_),
    .A2(_2900_),
    .A3(_1579_),
    .B1(_2897_),
    .X(_2975_));
 sky130_fd_sc_hd__a31o_1 _6344_ (.A1(_0743_),
    .A2(_2973_),
    .A3(_2974_),
    .B1(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__o21a_1 _6345_ (.A1(\core_0.execute.alu_mul_div.mul_res[8] ),
    .A2(_2952_),
    .B1(_2976_),
    .X(_0411_));
 sky130_fd_sc_hd__inv_2 _6346_ (.A(\core_0.execute.alu_mul_div.mul_res[9] ),
    .Y(_2977_));
 sky130_fd_sc_hd__mux4_1 _6347_ (.A0(_1550_),
    .A1(_1571_),
    .A2(_1579_),
    .A3(_1654_),
    .S0(_1206_),
    .S1(_1205_),
    .X(_2978_));
 sky130_fd_sc_hd__nand2_1 _6348_ (.A(_1204_),
    .B(_2978_),
    .Y(_2979_));
 sky130_fd_sc_hd__o211a_1 _6349_ (.A1(_1204_),
    .A2(_2936_),
    .B1(_2979_),
    .C1(_1803_),
    .X(_2980_));
 sky130_fd_sc_hd__o21bai_2 _6350_ (.A1(_1803_),
    .A2(_2902_),
    .B1_N(_2980_),
    .Y(_2981_));
 sky130_fd_sc_hd__nor2_1 _6351_ (.A(_2977_),
    .B(_2981_),
    .Y(_2982_));
 sky130_fd_sc_hd__nand2_1 _6352_ (.A(_2977_),
    .B(_2981_),
    .Y(_2983_));
 sky130_fd_sc_hd__and2b_1 _6353_ (.A_N(_2982_),
    .B(_2983_),
    .X(_2984_));
 sky130_fd_sc_hd__a21o_1 _6354_ (.A1(_2971_),
    .A2(_2972_),
    .B1(_2969_),
    .X(_2985_));
 sky130_fd_sc_hd__nand2_1 _6355_ (.A(_2984_),
    .B(_2985_),
    .Y(_2986_));
 sky130_fd_sc_hd__o21a_1 _6356_ (.A1(_2984_),
    .A2(_2985_),
    .B1(_0743_),
    .X(_2987_));
 sky130_fd_sc_hd__a32o_1 _6357_ (.A1(_2874_),
    .A2(_2002_),
    .A3(_1550_),
    .B1(_2986_),
    .B2(_2987_),
    .X(_2988_));
 sky130_fd_sc_hd__mux2_1 _6358_ (.A0(\core_0.execute.alu_mul_div.mul_res[9] ),
    .A1(_2988_),
    .S(_2952_),
    .X(_2989_));
 sky130_fd_sc_hd__clkbuf_1 _6359_ (.A(_2989_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_1 _6360_ (.A(_1435_),
    .B(_1581_),
    .Y(_2990_));
 sky130_fd_sc_hd__a211oi_1 _6361_ (.A1(_1435_),
    .A2(_1679_),
    .B1(_2990_),
    .C1(_1201_),
    .Y(_2991_));
 sky130_fd_sc_hd__a31o_1 _6362_ (.A1(_1202_),
    .A2(_1204_),
    .A3(_1646_),
    .B1(_2991_),
    .X(_2992_));
 sky130_fd_sc_hd__and2_1 _6363_ (.A(\core_0.execute.alu_mul_div.mul_res[10] ),
    .B(_2992_),
    .X(_2993_));
 sky130_fd_sc_hd__nor2_1 _6364_ (.A(\core_0.execute.alu_mul_div.mul_res[10] ),
    .B(_2992_),
    .Y(_2994_));
 sky130_fd_sc_hd__nor2_1 _6365_ (.A(_2993_),
    .B(_2994_),
    .Y(_2995_));
 sky130_fd_sc_hd__a21o_1 _6366_ (.A1(_2983_),
    .A2(_2985_),
    .B1(_2982_),
    .X(_2996_));
 sky130_fd_sc_hd__o21ai_1 _6367_ (.A1(_2995_),
    .A2(_2996_),
    .B1(_0743_),
    .Y(_2997_));
 sky130_fd_sc_hd__a21oi_1 _6368_ (.A1(_2995_),
    .A2(_2996_),
    .B1(_2997_),
    .Y(_2998_));
 sky130_fd_sc_hd__a31o_1 _6369_ (.A1(_2875_),
    .A2(_2900_),
    .A3(_1558_),
    .B1(_2898_),
    .X(_2999_));
 sky130_fd_sc_hd__o22a_1 _6370_ (.A1(\core_0.execute.alu_mul_div.mul_res[10] ),
    .A2(_2952_),
    .B1(_2998_),
    .B2(_2999_),
    .X(_0413_));
 sky130_fd_sc_hd__a21oi_1 _6371_ (.A1(_2995_),
    .A2(_2996_),
    .B1(_2993_),
    .Y(_3000_));
 sky130_fd_sc_hd__mux4_1 _6372_ (.A0(_1558_),
    .A1(_1594_),
    .A2(_1579_),
    .A3(_1550_),
    .S0(_1560_),
    .S1(_1206_),
    .X(_3001_));
 sky130_fd_sc_hd__nor2_1 _6373_ (.A(_1435_),
    .B(_3001_),
    .Y(_3002_));
 sky130_fd_sc_hd__a211o_1 _6374_ (.A1(_1435_),
    .A2(_2954_),
    .B1(_3002_),
    .C1(_1202_),
    .X(_3003_));
 sky130_fd_sc_hd__o21ai_1 _6375_ (.A1(_1803_),
    .A2(_2928_),
    .B1(_3003_),
    .Y(_3004_));
 sky130_fd_sc_hd__and2_1 _6376_ (.A(\core_0.execute.alu_mul_div.mul_res[11] ),
    .B(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__or2_1 _6377_ (.A(\core_0.execute.alu_mul_div.mul_res[11] ),
    .B(_3004_),
    .X(_3006_));
 sky130_fd_sc_hd__inv_2 _6378_ (.A(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__or3_1 _6379_ (.A(_3000_),
    .B(_3005_),
    .C(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__o21ai_1 _6380_ (.A1(_3005_),
    .A2(_3007_),
    .B1(_3000_),
    .Y(_3009_));
 sky130_fd_sc_hd__a32o_1 _6381_ (.A1(_2875_),
    .A2(_2900_),
    .A3(_1594_),
    .B1(_2898_),
    .B2(\core_0.execute.alu_mul_div.mul_res[11] ),
    .X(_3010_));
 sky130_fd_sc_hd__a31o_1 _6382_ (.A1(_2892_),
    .A2(_3008_),
    .A3(_3009_),
    .B1(_3010_),
    .X(_0414_));
 sky130_fd_sc_hd__inv_2 _6383_ (.A(_2924_),
    .Y(_3011_));
 sky130_fd_sc_hd__mux4_1 _6384_ (.A0(_1580_),
    .A1(_1662_),
    .A2(_1595_),
    .A3(_1561_),
    .S0(_1207_),
    .S1(_1204_),
    .X(_3012_));
 sky130_fd_sc_hd__mux2_1 _6385_ (.A0(_3011_),
    .A1(_3012_),
    .S(_1803_),
    .X(_3013_));
 sky130_fd_sc_hd__and2_1 _6386_ (.A(\core_0.execute.alu_mul_div.mul_res[12] ),
    .B(_3013_),
    .X(_3014_));
 sky130_fd_sc_hd__nor2_1 _6387_ (.A(\core_0.execute.alu_mul_div.mul_res[12] ),
    .B(_3013_),
    .Y(_3015_));
 sky130_fd_sc_hd__nor2_1 _6388_ (.A(_3014_),
    .B(_3015_),
    .Y(_3016_));
 sky130_fd_sc_hd__a211o_1 _6389_ (.A1(_2995_),
    .A2(_2996_),
    .B1(_3005_),
    .C1(_2993_),
    .X(_3017_));
 sky130_fd_sc_hd__nand2_1 _6390_ (.A(_3006_),
    .B(_3017_),
    .Y(_3018_));
 sky130_fd_sc_hd__xnor2_1 _6391_ (.A(_3016_),
    .B(_3018_),
    .Y(_3019_));
 sky130_fd_sc_hd__a31o_1 _6392_ (.A1(_2874_),
    .A2(_2900_),
    .A3(_1588_),
    .B1(_2897_),
    .X(_3020_));
 sky130_fd_sc_hd__a21o_1 _6393_ (.A1(_0743_),
    .A2(_3019_),
    .B1(_3020_),
    .X(_3021_));
 sky130_fd_sc_hd__o21a_1 _6394_ (.A1(\core_0.execute.alu_mul_div.mul_res[12] ),
    .A2(_2952_),
    .B1(_3021_),
    .X(_0415_));
 sky130_fd_sc_hd__and3_1 _6395_ (.A(_3006_),
    .B(_3016_),
    .C(_3017_),
    .X(_3022_));
 sky130_fd_sc_hd__inv_2 _6396_ (.A(\core_0.execute.alu_mul_div.mul_res[13] ),
    .Y(_3023_));
 sky130_fd_sc_hd__mux4_1 _6397_ (.A0(_1756_),
    .A1(_1757_),
    .A2(_1920_),
    .A3(_1914_),
    .S0(_1560_),
    .S1(_1207_),
    .X(_3024_));
 sky130_fd_sc_hd__nand2_1 _6398_ (.A(_1435_),
    .B(_2978_),
    .Y(_3025_));
 sky130_fd_sc_hd__o211a_1 _6399_ (.A1(_1435_),
    .A2(_3024_),
    .B1(_3025_),
    .C1(_1803_),
    .X(_3026_));
 sky130_fd_sc_hd__a21o_1 _6400_ (.A1(_1202_),
    .A2(_2938_),
    .B1(_3026_),
    .X(_3027_));
 sky130_fd_sc_hd__or2_1 _6401_ (.A(_3023_),
    .B(_3027_),
    .X(_3028_));
 sky130_fd_sc_hd__nand2_1 _6402_ (.A(_3023_),
    .B(_3027_),
    .Y(_3029_));
 sky130_fd_sc_hd__nand2_1 _6403_ (.A(_3028_),
    .B(_3029_),
    .Y(_3030_));
 sky130_fd_sc_hd__o21bai_1 _6404_ (.A1(_3014_),
    .A2(_3022_),
    .B1_N(_3030_),
    .Y(_3031_));
 sky130_fd_sc_hd__or3b_1 _6405_ (.A(_3014_),
    .B(_3022_),
    .C_N(_3030_),
    .X(_3032_));
 sky130_fd_sc_hd__and3_1 _6406_ (.A(_2874_),
    .B(_2002_),
    .C(_1601_),
    .X(_3033_));
 sky130_fd_sc_hd__a31o_1 _6407_ (.A1(_0743_),
    .A2(_3031_),
    .A3(_3032_),
    .B1(_3033_),
    .X(_3034_));
 sky130_fd_sc_hd__mux2_1 _6408_ (.A0(\core_0.execute.alu_mul_div.mul_res[13] ),
    .A1(_3034_),
    .S(_2952_),
    .X(_3035_));
 sky130_fd_sc_hd__clkbuf_1 _6409_ (.A(_3035_),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _6410_ (.A(\core_0.execute.alu_mul_div.mul_res[14] ),
    .B(_1682_),
    .X(_3036_));
 sky130_fd_sc_hd__nor2_1 _6411_ (.A(\core_0.execute.alu_mul_div.mul_res[14] ),
    .B(_1682_),
    .Y(_3037_));
 sky130_fd_sc_hd__or2_1 _6412_ (.A(_3036_),
    .B(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__a21oi_1 _6413_ (.A1(_3028_),
    .A2(_3031_),
    .B1(_3038_),
    .Y(_3039_));
 sky130_fd_sc_hd__a31o_1 _6414_ (.A1(_3028_),
    .A2(_3031_),
    .A3(_3038_),
    .B1(_2874_),
    .X(_3040_));
 sky130_fd_sc_hd__nor2_1 _6415_ (.A(_3039_),
    .B(_3040_),
    .Y(_3041_));
 sky130_fd_sc_hd__a31o_1 _6416_ (.A1(_2875_),
    .A2(_2900_),
    .A3(_1841_),
    .B1(_2898_),
    .X(_3042_));
 sky130_fd_sc_hd__o22a_1 _6417_ (.A1(\core_0.execute.alu_mul_div.mul_res[14] ),
    .A2(_2952_),
    .B1(_3041_),
    .B2(_3042_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _6418_ (.A0(_1588_),
    .A1(_1601_),
    .S(_1560_),
    .X(_3043_));
 sky130_fd_sc_hd__a21o_1 _6419_ (.A1(_1207_),
    .A2(_3043_),
    .B1(_1435_),
    .X(_3044_));
 sky130_fd_sc_hd__a221o_1 _6420_ (.A1(_1797_),
    .A2(_1542_),
    .B1(_1602_),
    .B2(_1841_),
    .C1(_3044_),
    .X(_3045_));
 sky130_fd_sc_hd__o21ai_1 _6421_ (.A1(_1799_),
    .A2(_3001_),
    .B1(_3045_),
    .Y(_3046_));
 sky130_fd_sc_hd__mux2_1 _6422_ (.A0(_2955_),
    .A1(_3046_),
    .S(_1803_),
    .X(_3047_));
 sky130_fd_sc_hd__xnor2_1 _6423_ (.A(\core_0.execute.alu_mul_div.mul_res[15] ),
    .B(_3047_),
    .Y(_3048_));
 sky130_fd_sc_hd__or3_1 _6424_ (.A(_3036_),
    .B(_3039_),
    .C(_3048_),
    .X(_3049_));
 sky130_fd_sc_hd__o21ai_1 _6425_ (.A1(_3036_),
    .A2(_3039_),
    .B1(_3048_),
    .Y(_3050_));
 sky130_fd_sc_hd__a32o_1 _6426_ (.A1(_2875_),
    .A2(_2900_),
    .A3(_1542_),
    .B1(_2898_),
    .B2(\core_0.execute.alu_mul_div.mul_res[15] ),
    .X(_3051_));
 sky130_fd_sc_hd__a31o_1 _6427_ (.A1(_2892_),
    .A2(_3049_),
    .A3(_3050_),
    .B1(_3051_),
    .X(_0418_));
 sky130_fd_sc_hd__nor2_1 _6428_ (.A(_1128_),
    .B(_0740_),
    .Y(_0419_));
 sky130_fd_sc_hd__nor2_1 _6429_ (.A(_1210_),
    .B(_1516_),
    .Y(_3052_));
 sky130_fd_sc_hd__o21a_1 _6430_ (.A1(\core_0.execute.alu_mul_div.div_res[0] ),
    .A2(_3052_),
    .B1(_1430_),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_2 _6431_ (.A(_1803_),
    .B(_1516_),
    .Y(_3053_));
 sky130_fd_sc_hd__a31o_1 _6432_ (.A1(_1436_),
    .A2(_1645_),
    .A3(_3053_),
    .B1(\core_0.execute.alu_mul_div.div_res[1] ),
    .X(_3054_));
 sky130_fd_sc_hd__and2_1 _6433_ (.A(_1474_),
    .B(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__clkbuf_1 _6434_ (.A(_3055_),
    .X(_0421_));
 sky130_fd_sc_hd__buf_2 _6435_ (.A(_0742_),
    .X(_3056_));
 sky130_fd_sc_hd__a31o_1 _6436_ (.A1(_1436_),
    .A2(_1602_),
    .A3(_3053_),
    .B1(\core_0.execute.alu_mul_div.div_res[2] ),
    .X(_3057_));
 sky130_fd_sc_hd__and2_1 _6437_ (.A(_3056_),
    .B(_3057_),
    .X(_3058_));
 sky130_fd_sc_hd__clkbuf_1 _6438_ (.A(_3058_),
    .X(_0422_));
 sky130_fd_sc_hd__a31o_1 _6439_ (.A1(_1436_),
    .A2(_1797_),
    .A3(_3053_),
    .B1(\core_0.execute.alu_mul_div.div_res[3] ),
    .X(_3059_));
 sky130_fd_sc_hd__and2_1 _6440_ (.A(_3056_),
    .B(_3059_),
    .X(_3060_));
 sky130_fd_sc_hd__clkbuf_1 _6441_ (.A(_3060_),
    .X(_0423_));
 sky130_fd_sc_hd__and3_1 _6442_ (.A(_1799_),
    .B(_1437_),
    .C(_3053_),
    .X(_3061_));
 sky130_fd_sc_hd__o21a_1 _6443_ (.A1(\core_0.execute.alu_mul_div.div_res[4] ),
    .A2(_3061_),
    .B1(_1430_),
    .X(_0424_));
 sky130_fd_sc_hd__a31o_1 _6444_ (.A1(_1799_),
    .A2(_1645_),
    .A3(_3053_),
    .B1(\core_0.execute.alu_mul_div.div_res[5] ),
    .X(_3062_));
 sky130_fd_sc_hd__and2_1 _6445_ (.A(_3056_),
    .B(_3062_),
    .X(_3063_));
 sky130_fd_sc_hd__clkbuf_1 _6446_ (.A(_3063_),
    .X(_0425_));
 sky130_fd_sc_hd__a31o_1 _6447_ (.A1(_1799_),
    .A2(_1602_),
    .A3(_3053_),
    .B1(\core_0.execute.alu_mul_div.div_res[6] ),
    .X(_3064_));
 sky130_fd_sc_hd__and2_1 _6448_ (.A(_3056_),
    .B(_3064_),
    .X(_3065_));
 sky130_fd_sc_hd__clkbuf_1 _6449_ (.A(_3065_),
    .X(_0426_));
 sky130_fd_sc_hd__and2_1 _6450_ (.A(_1409_),
    .B(_1412_),
    .X(_3066_));
 sky130_fd_sc_hd__and4_1 _6451_ (.A(_1202_),
    .B(_1799_),
    .C(_1797_),
    .D(_3066_),
    .X(_3067_));
 sky130_fd_sc_hd__o21a_1 _6452_ (.A1(\core_0.execute.alu_mul_div.div_res[7] ),
    .A2(_3067_),
    .B1(_1430_),
    .X(_0427_));
 sky130_fd_sc_hd__a31o_1 _6453_ (.A1(_1803_),
    .A2(_1209_),
    .A3(_3066_),
    .B1(\core_0.execute.alu_mul_div.div_res[8] ),
    .X(_3068_));
 sky130_fd_sc_hd__and2_1 _6454_ (.A(_3056_),
    .B(_3068_),
    .X(_3069_));
 sky130_fd_sc_hd__clkbuf_1 _6455_ (.A(_3069_),
    .X(_0428_));
 sky130_fd_sc_hd__nor2_4 _6456_ (.A(_1202_),
    .B(_1516_),
    .Y(_3070_));
 sky130_fd_sc_hd__a31o_1 _6457_ (.A1(_1436_),
    .A2(_1645_),
    .A3(_3070_),
    .B1(\core_0.execute.alu_mul_div.div_res[9] ),
    .X(_3071_));
 sky130_fd_sc_hd__and2_1 _6458_ (.A(_3056_),
    .B(_3071_),
    .X(_3072_));
 sky130_fd_sc_hd__clkbuf_1 _6459_ (.A(_3072_),
    .X(_0429_));
 sky130_fd_sc_hd__a31o_1 _6460_ (.A1(_1436_),
    .A2(_1602_),
    .A3(_3070_),
    .B1(\core_0.execute.alu_mul_div.div_res[10] ),
    .X(_3073_));
 sky130_fd_sc_hd__and2_1 _6461_ (.A(_3056_),
    .B(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__clkbuf_1 _6462_ (.A(_3074_),
    .X(_0430_));
 sky130_fd_sc_hd__a31o_1 _6463_ (.A1(_1436_),
    .A2(_1797_),
    .A3(_3070_),
    .B1(\core_0.execute.alu_mul_div.div_res[11] ),
    .X(_3075_));
 sky130_fd_sc_hd__and2_1 _6464_ (.A(_3056_),
    .B(_3075_),
    .X(_3076_));
 sky130_fd_sc_hd__clkbuf_1 _6465_ (.A(_3076_),
    .X(_0431_));
 sky130_fd_sc_hd__and3_1 _6466_ (.A(_1799_),
    .B(_1437_),
    .C(_3070_),
    .X(_3077_));
 sky130_fd_sc_hd__o21a_1 _6467_ (.A1(\core_0.execute.alu_mul_div.div_res[12] ),
    .A2(_3077_),
    .B1(_1430_),
    .X(_0432_));
 sky130_fd_sc_hd__a31o_1 _6468_ (.A1(_1799_),
    .A2(_1645_),
    .A3(_3070_),
    .B1(\core_0.execute.alu_mul_div.div_res[13] ),
    .X(_3078_));
 sky130_fd_sc_hd__and2_1 _6469_ (.A(_3056_),
    .B(_3078_),
    .X(_3079_));
 sky130_fd_sc_hd__clkbuf_1 _6470_ (.A(_3079_),
    .X(_0433_));
 sky130_fd_sc_hd__a31o_1 _6471_ (.A1(_1799_),
    .A2(_1602_),
    .A3(_3070_),
    .B1(\core_0.execute.alu_mul_div.div_res[14] ),
    .X(_3080_));
 sky130_fd_sc_hd__and2_1 _6472_ (.A(_3056_),
    .B(_3080_),
    .X(_3081_));
 sky130_fd_sc_hd__clkbuf_1 _6473_ (.A(_3081_),
    .X(_0434_));
 sky130_fd_sc_hd__a31o_1 _6474_ (.A1(_1799_),
    .A2(_1797_),
    .A3(_3070_),
    .B1(\core_0.execute.alu_mul_div.div_res[15] ),
    .X(_3082_));
 sky130_fd_sc_hd__and2_1 _6475_ (.A(_0742_),
    .B(_3082_),
    .X(_3083_));
 sky130_fd_sc_hd__clkbuf_1 _6476_ (.A(_3083_),
    .X(_0435_));
 sky130_fd_sc_hd__o21ai_1 _6477_ (.A1(net79),
    .A2(_1693_),
    .B1(_1691_),
    .Y(_3084_));
 sky130_fd_sc_hd__a21o_1 _6478_ (.A1(net79),
    .A2(_1693_),
    .B1(_3084_),
    .X(_3085_));
 sky130_fd_sc_hd__nor2_2 _6479_ (.A(_1038_),
    .B(_1152_),
    .Y(_3086_));
 sky130_fd_sc_hd__buf_2 _6480_ (.A(_3086_),
    .X(_3087_));
 sky130_fd_sc_hd__and2_1 _6481_ (.A(_1789_),
    .B(_1152_),
    .X(_3088_));
 sky130_fd_sc_hd__clkbuf_4 _6482_ (.A(_3088_),
    .X(_3089_));
 sky130_fd_sc_hd__a221o_1 _6483_ (.A1(\core_0.execute.sreg_irq_pc.o_d[1] ),
    .A2(_1154_),
    .B1(net201),
    .B2(_3089_),
    .C1(_1691_),
    .X(_3090_));
 sky130_fd_sc_hd__a21o_1 _6484_ (.A1(_3087_),
    .A2(_2138_),
    .B1(_3090_),
    .X(_3091_));
 sky130_fd_sc_hd__and3_1 _6485_ (.A(_2870_),
    .B(_3085_),
    .C(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__clkbuf_1 _6486_ (.A(_3092_),
    .X(_0436_));
 sky130_fd_sc_hd__a21oi_1 _6487_ (.A1(net79),
    .A2(net72),
    .B1(net80),
    .Y(_3093_));
 sky130_fd_sc_hd__and3_1 _6488_ (.A(net80),
    .B(net79),
    .C(net72),
    .X(_3094_));
 sky130_fd_sc_hd__or3b_4 _6489_ (.A(_1685_),
    .B(_1690_),
    .C_N(_1027_),
    .X(_3095_));
 sky130_fd_sc_hd__or3_1 _6490_ (.A(_3093_),
    .B(_3094_),
    .C(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__o31ai_4 _6491_ (.A1(\core_0.dec_jump_cond_code[4] ),
    .A2(\core_0.dec_pc_inc ),
    .A3(_1039_),
    .B1(_1071_),
    .Y(_3097_));
 sky130_fd_sc_hd__a22o_1 _6492_ (.A1(\core_0.execute.sreg_irq_pc.o_d[2] ),
    .A2(_1154_),
    .B1(net202),
    .B2(_3089_),
    .X(_3098_));
 sky130_fd_sc_hd__a21oi_1 _6493_ (.A1(_3087_),
    .A2(_2187_),
    .B1(_3098_),
    .Y(_3099_));
 sky130_fd_sc_hd__o2bb2a_1 _6494_ (.A1_N(net80),
    .A2_N(_3097_),
    .B1(_3099_),
    .B2(_1692_),
    .X(_3100_));
 sky130_fd_sc_hd__a21oi_1 _6495_ (.A1(_3096_),
    .A2(_3100_),
    .B1(_1168_),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2_1 _6496_ (.A(_1687_),
    .B(_3094_),
    .Y(_3101_));
 sky130_fd_sc_hd__xor2_1 _6497_ (.A(net81),
    .B(_3101_),
    .X(_3102_));
 sky130_fd_sc_hd__nand2_1 _6498_ (.A(_1692_),
    .B(_3102_),
    .Y(_3103_));
 sky130_fd_sc_hd__a21o_1 _6499_ (.A1(net203),
    .A2(_3089_),
    .B1(_2205_),
    .X(_3104_));
 sky130_fd_sc_hd__a211o_1 _6500_ (.A1(_3087_),
    .A2(_2241_),
    .B1(_3104_),
    .C1(_1791_),
    .X(_3105_));
 sky130_fd_sc_hd__and3_1 _6501_ (.A(_2870_),
    .B(_3103_),
    .C(_3105_),
    .X(_3106_));
 sky130_fd_sc_hd__clkbuf_1 _6502_ (.A(_3106_),
    .X(_0438_));
 sky130_fd_sc_hd__a21oi_1 _6503_ (.A1(net81),
    .A2(_3094_),
    .B1(net82),
    .Y(_3107_));
 sky130_fd_sc_hd__and3_1 _6504_ (.A(net82),
    .B(net81),
    .C(_3094_),
    .X(_3108_));
 sky130_fd_sc_hd__or3_1 _6505_ (.A(_3095_),
    .B(_3107_),
    .C(_3108_),
    .X(_3109_));
 sky130_fd_sc_hd__nand2_1 _6506_ (.A(_3086_),
    .B(_2266_),
    .Y(_3110_));
 sky130_fd_sc_hd__o211a_1 _6507_ (.A1(_0633_),
    .A2(_1790_),
    .B1(_2273_),
    .C1(_3110_),
    .X(_3111_));
 sky130_fd_sc_hd__o2bb2a_1 _6508_ (.A1_N(net82),
    .A2_N(_3097_),
    .B1(_3111_),
    .B2(_1692_),
    .X(_3112_));
 sky130_fd_sc_hd__a21oi_1 _6509_ (.A1(_3109_),
    .A2(_3112_),
    .B1(_1168_),
    .Y(_0439_));
 sky130_fd_sc_hd__nand2_1 _6510_ (.A(_1687_),
    .B(_3108_),
    .Y(_3113_));
 sky130_fd_sc_hd__xnor2_1 _6511_ (.A(_1813_),
    .B(_3113_),
    .Y(_3114_));
 sky130_fd_sc_hd__nand2_1 _6512_ (.A(_1692_),
    .B(_3114_),
    .Y(_3115_));
 sky130_fd_sc_hd__a22o_1 _6513_ (.A1(\core_0.execute.sreg_irq_pc.o_d[5] ),
    .A2(_1038_),
    .B1(net205),
    .B2(_3088_),
    .X(_3116_));
 sky130_fd_sc_hd__a211o_1 _6514_ (.A1(_3087_),
    .A2(_2298_),
    .B1(_3116_),
    .C1(_1791_),
    .X(_3117_));
 sky130_fd_sc_hd__and3_1 _6515_ (.A(_2870_),
    .B(_3115_),
    .C(_3117_),
    .X(_3118_));
 sky130_fd_sc_hd__clkbuf_1 _6516_ (.A(_3118_),
    .X(_0440_));
 sky130_fd_sc_hd__and3_1 _6517_ (.A(net84),
    .B(net83),
    .C(_3108_),
    .X(_3119_));
 sky130_fd_sc_hd__a21oi_1 _6518_ (.A1(net83),
    .A2(_3108_),
    .B1(net84),
    .Y(_3120_));
 sky130_fd_sc_hd__or3_1 _6519_ (.A(_3095_),
    .B(_3119_),
    .C(_3120_),
    .X(_3121_));
 sky130_fd_sc_hd__a22o_1 _6520_ (.A1(\core_0.execute.sreg_irq_pc.o_d[6] ),
    .A2(_1154_),
    .B1(net206),
    .B2(_3089_),
    .X(_3122_));
 sky130_fd_sc_hd__a21oi_1 _6521_ (.A1(_3087_),
    .A2(_2341_),
    .B1(_3122_),
    .Y(_3123_));
 sky130_fd_sc_hd__o2bb2a_1 _6522_ (.A1_N(net84),
    .A2_N(_3097_),
    .B1(_3123_),
    .B2(_1791_),
    .X(_3124_));
 sky130_fd_sc_hd__a21oi_1 _6523_ (.A1(_3121_),
    .A2(_3124_),
    .B1(_1168_),
    .Y(_0441_));
 sky130_fd_sc_hd__nand2_1 _6524_ (.A(_1687_),
    .B(_3119_),
    .Y(_3125_));
 sky130_fd_sc_hd__xnor2_1 _6525_ (.A(_1819_),
    .B(_3125_),
    .Y(_3126_));
 sky130_fd_sc_hd__nand2_1 _6526_ (.A(_1692_),
    .B(_3126_),
    .Y(_3127_));
 sky130_fd_sc_hd__a22o_1 _6527_ (.A1(\core_0.execute.sreg_irq_pc.o_d[7] ),
    .A2(_1038_),
    .B1(net207),
    .B2(_3088_),
    .X(_3128_));
 sky130_fd_sc_hd__a211o_1 _6528_ (.A1(_3087_),
    .A2(_2367_),
    .B1(_3128_),
    .C1(_1791_),
    .X(_3129_));
 sky130_fd_sc_hd__and3_1 _6529_ (.A(_2869_),
    .B(_3127_),
    .C(_3129_),
    .X(_3130_));
 sky130_fd_sc_hd__clkbuf_1 _6530_ (.A(_3130_),
    .X(_0442_));
 sky130_fd_sc_hd__and3_1 _6531_ (.A(net86),
    .B(net85),
    .C(_3119_),
    .X(_3131_));
 sky130_fd_sc_hd__a21oi_1 _6532_ (.A1(net85),
    .A2(_3119_),
    .B1(net86),
    .Y(_3132_));
 sky130_fd_sc_hd__or3_1 _6533_ (.A(_3095_),
    .B(_3131_),
    .C(_3132_),
    .X(_3133_));
 sky130_fd_sc_hd__a22o_1 _6534_ (.A1(\core_0.execute.sreg_irq_pc.o_d[8] ),
    .A2(_1154_),
    .B1(net208),
    .B2(_3089_),
    .X(_3134_));
 sky130_fd_sc_hd__a21oi_1 _6535_ (.A1(_3087_),
    .A2(_2396_),
    .B1(_3134_),
    .Y(_3135_));
 sky130_fd_sc_hd__o2bb2a_1 _6536_ (.A1_N(net86),
    .A2_N(_3097_),
    .B1(_3135_),
    .B2(_1791_),
    .X(_3136_));
 sky130_fd_sc_hd__a21oi_1 _6537_ (.A1(_3133_),
    .A2(_3136_),
    .B1(_1168_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand2_1 _6538_ (.A(_1687_),
    .B(_3131_),
    .Y(_3137_));
 sky130_fd_sc_hd__xor2_1 _6539_ (.A(net87),
    .B(_3137_),
    .X(_3138_));
 sky130_fd_sc_hd__nand2_1 _6540_ (.A(_1692_),
    .B(_3138_),
    .Y(_3139_));
 sky130_fd_sc_hd__a21o_1 _6541_ (.A1(net209),
    .A2(_3089_),
    .B1(_2433_),
    .X(_3140_));
 sky130_fd_sc_hd__a211o_1 _6542_ (.A1(_3087_),
    .A2(_2427_),
    .B1(_3140_),
    .C1(_1691_),
    .X(_3141_));
 sky130_fd_sc_hd__and3_1 _6543_ (.A(_2869_),
    .B(_3139_),
    .C(_3141_),
    .X(_3142_));
 sky130_fd_sc_hd__clkbuf_1 _6544_ (.A(_3142_),
    .X(_0444_));
 sky130_fd_sc_hd__and3_1 _6545_ (.A(net73),
    .B(net87),
    .C(_3131_),
    .X(_3143_));
 sky130_fd_sc_hd__a21oi_1 _6546_ (.A1(net87),
    .A2(_3131_),
    .B1(net73),
    .Y(_3144_));
 sky130_fd_sc_hd__or3_1 _6547_ (.A(_3095_),
    .B(_3143_),
    .C(_3144_),
    .X(_3145_));
 sky130_fd_sc_hd__nand2_1 _6548_ (.A(_3086_),
    .B(_2459_),
    .Y(_3146_));
 sky130_fd_sc_hd__o211a_1 _6549_ (.A1(_0592_),
    .A2(_1790_),
    .B1(_2464_),
    .C1(_3146_),
    .X(_3147_));
 sky130_fd_sc_hd__o2bb2a_1 _6550_ (.A1_N(net73),
    .A2_N(_3097_),
    .B1(_3147_),
    .B2(_1791_),
    .X(_3148_));
 sky130_fd_sc_hd__a21oi_1 _6551_ (.A1(_3145_),
    .A2(_3148_),
    .B1(_1168_),
    .Y(_0445_));
 sky130_fd_sc_hd__o221a_1 _6552_ (.A1(_1340_),
    .A2(_1790_),
    .B1(_2494_),
    .B2(_1695_),
    .C1(_2499_),
    .X(_3149_));
 sky130_fd_sc_hd__nand2_1 _6553_ (.A(_1687_),
    .B(_3143_),
    .Y(_3150_));
 sky130_fd_sc_hd__xnor2_1 _6554_ (.A(_1825_),
    .B(_3150_),
    .Y(_3151_));
 sky130_fd_sc_hd__mux2_1 _6555_ (.A0(_3149_),
    .A1(_3151_),
    .S(_1791_),
    .X(_3152_));
 sky130_fd_sc_hd__nor2_1 _6556_ (.A(_1168_),
    .B(_3152_),
    .Y(_0446_));
 sky130_fd_sc_hd__and3_1 _6557_ (.A(net75),
    .B(net74),
    .C(_3143_),
    .X(_3153_));
 sky130_fd_sc_hd__a21oi_1 _6558_ (.A1(net74),
    .A2(_3143_),
    .B1(net75),
    .Y(_3154_));
 sky130_fd_sc_hd__or3_1 _6559_ (.A(_3095_),
    .B(_3153_),
    .C(_3154_),
    .X(_3155_));
 sky130_fd_sc_hd__a221oi_2 _6560_ (.A1(net197),
    .A2(_3089_),
    .B1(_2523_),
    .B2(_3086_),
    .C1(_2529_),
    .Y(_3156_));
 sky130_fd_sc_hd__o2bb2a_1 _6561_ (.A1_N(net75),
    .A2_N(_3097_),
    .B1(_3156_),
    .B2(_1791_),
    .X(_3157_));
 sky130_fd_sc_hd__a21oi_1 _6562_ (.A1(_3155_),
    .A2(_3157_),
    .B1(_1168_),
    .Y(_0447_));
 sky130_fd_sc_hd__nor2_1 _6563_ (.A(_1695_),
    .B(_2562_),
    .Y(_3158_));
 sky130_fd_sc_hd__a221o_1 _6564_ (.A1(\core_0.execute.sreg_irq_pc.o_d[13] ),
    .A2(_1154_),
    .B1(net198),
    .B2(_3089_),
    .C1(_1692_),
    .X(_3159_));
 sky130_fd_sc_hd__nand2_1 _6565_ (.A(_1687_),
    .B(_3153_),
    .Y(_3160_));
 sky130_fd_sc_hd__xnor2_1 _6566_ (.A(_1828_),
    .B(_3160_),
    .Y(_3161_));
 sky130_fd_sc_hd__nand2_1 _6567_ (.A(_1692_),
    .B(_3161_),
    .Y(_3162_));
 sky130_fd_sc_hd__o211a_1 _6568_ (.A1(_3158_),
    .A2(_3159_),
    .B1(_3162_),
    .C1(_2870_),
    .X(_0448_));
 sky130_fd_sc_hd__and3_1 _6569_ (.A(net77),
    .B(net76),
    .C(_3153_),
    .X(_3163_));
 sky130_fd_sc_hd__a21oi_1 _6570_ (.A1(net76),
    .A2(_3153_),
    .B1(net77),
    .Y(_3164_));
 sky130_fd_sc_hd__or3_1 _6571_ (.A(_3095_),
    .B(_3163_),
    .C(_3164_),
    .X(_3165_));
 sky130_fd_sc_hd__a22o_1 _6572_ (.A1(\core_0.execute.sreg_irq_pc.o_d[14] ),
    .A2(_1154_),
    .B1(net199),
    .B2(_3089_),
    .X(_3166_));
 sky130_fd_sc_hd__a21oi_1 _6573_ (.A1(_3087_),
    .A2(_2585_),
    .B1(_3166_),
    .Y(_3167_));
 sky130_fd_sc_hd__o2bb2a_1 _6574_ (.A1_N(net77),
    .A2_N(_3097_),
    .B1(_3167_),
    .B2(_1791_),
    .X(_3168_));
 sky130_fd_sc_hd__a21oi_1 _6575_ (.A1(_3165_),
    .A2(_3168_),
    .B1(_1168_),
    .Y(_0449_));
 sky130_fd_sc_hd__xnor2_1 _6576_ (.A(net78),
    .B(_3163_),
    .Y(_3169_));
 sky130_fd_sc_hd__a221o_1 _6577_ (.A1(\core_0.execute.sreg_irq_pc.o_d[15] ),
    .A2(_1154_),
    .B1(net200),
    .B2(_3089_),
    .C1(_1691_),
    .X(_3170_));
 sky130_fd_sc_hd__a21oi_1 _6578_ (.A1(_3087_),
    .A2(_2615_),
    .B1(_3170_),
    .Y(_3171_));
 sky130_fd_sc_hd__a21oi_1 _6579_ (.A1(_1692_),
    .A2(_3169_),
    .B1(_3171_),
    .Y(_3172_));
 sky130_fd_sc_hd__or2b_1 _6580_ (.A(net78),
    .B_N(_3097_),
    .X(_3173_));
 sky130_fd_sc_hd__o211a_1 _6581_ (.A1(_3097_),
    .A2(_3172_),
    .B1(_3173_),
    .C1(_2870_),
    .X(_0450_));
 sky130_fd_sc_hd__and2_1 _6582_ (.A(\core_0.dec_sreg_store ),
    .B(_2079_),
    .X(_3174_));
 sky130_fd_sc_hd__clkbuf_4 _6583_ (.A(_3174_),
    .X(_3175_));
 sky130_fd_sc_hd__o21a_2 _6584_ (.A1(\core_0.dec_alu_flags_ie ),
    .A2(_3175_),
    .B1(_1027_),
    .X(_3176_));
 sky130_fd_sc_hd__or2_1 _6585_ (.A(_2582_),
    .B(_2611_),
    .X(_3177_));
 sky130_fd_sc_hd__nand2_1 _6586_ (.A(_2520_),
    .B(_2559_),
    .Y(_3178_));
 sky130_fd_sc_hd__nand3_1 _6587_ (.A(_2393_),
    .B(_2419_),
    .C(_2424_),
    .Y(_3179_));
 sky130_fd_sc_hd__and3_1 _6588_ (.A(_2184_),
    .B(_2225_),
    .C(_2237_),
    .X(_3180_));
 sky130_fd_sc_hd__or4b_1 _6589_ (.A(_1782_),
    .B(_2134_),
    .C(_3175_),
    .D_N(_3180_),
    .X(_3181_));
 sky130_fd_sc_hd__clkinv_2 _6590_ (.A(_2364_),
    .Y(_3182_));
 sky130_fd_sc_hd__and3b_1 _6591_ (.A_N(_2263_),
    .B(_2338_),
    .C(_3182_),
    .X(_3183_));
 sky130_fd_sc_hd__or4b_1 _6592_ (.A(_2295_),
    .B(_3179_),
    .C(_3181_),
    .D_N(_3183_),
    .X(_3184_));
 sky130_fd_sc_hd__or2_1 _6593_ (.A(_2456_),
    .B(_2491_),
    .X(_3185_));
 sky130_fd_sc_hd__or4_1 _6594_ (.A(_3177_),
    .B(_3178_),
    .C(_3184_),
    .D(_3185_),
    .X(_3186_));
 sky130_fd_sc_hd__nand2_1 _6595_ (.A(net194),
    .B(_3175_),
    .Y(_3187_));
 sky130_fd_sc_hd__a31o_1 _6596_ (.A1(_3186_),
    .A2(_3187_),
    .A3(_3176_),
    .B1(_1122_),
    .X(_3188_));
 sky130_fd_sc_hd__o21ba_1 _6597_ (.A1(\core_0.execute.alu_flag_reg.o_d[0] ),
    .A2(_3176_),
    .B1_N(_3188_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _6598_ (.A0(_2014_),
    .A1(_0655_),
    .S(_3175_),
    .X(_3189_));
 sky130_fd_sc_hd__nand2_1 _6599_ (.A(_3176_),
    .B(_3189_),
    .Y(_3190_));
 sky130_fd_sc_hd__o211a_1 _6600_ (.A1(\core_0.execute.alu_flag_reg.o_d[1] ),
    .A2(_3176_),
    .B1(_3190_),
    .C1(_2861_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _6601_ (.A0(_2611_),
    .A1(net202),
    .S(_3175_),
    .X(_3191_));
 sky130_fd_sc_hd__mux2_1 _6602_ (.A0(\core_0.execute.alu_flag_reg.o_d[2] ),
    .A1(_3191_),
    .S(_3176_),
    .X(_3192_));
 sky130_fd_sc_hd__and2_1 _6603_ (.A(_1190_),
    .B(_3192_),
    .X(_3193_));
 sky130_fd_sc_hd__clkbuf_1 _6604_ (.A(_3193_),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_1 _6605_ (.A(\core_0.execute.alu_flag_reg.o_d[3] ),
    .B(_3176_),
    .Y(_3194_));
 sky130_fd_sc_hd__a21oi_1 _6606_ (.A1(_0978_),
    .A2(_1934_),
    .B1(_3175_),
    .Y(_3195_));
 sky130_fd_sc_hd__o21ai_1 _6607_ (.A1(_0978_),
    .A2(_1934_),
    .B1(_3195_),
    .Y(_3196_));
 sky130_fd_sc_hd__a211o_1 _6608_ (.A1(_0978_),
    .A2(_2596_),
    .B1(_2610_),
    .C1(_1542_),
    .X(_3197_));
 sky130_fd_sc_hd__a21bo_1 _6609_ (.A1(_1542_),
    .A2(_2611_),
    .B1_N(_3197_),
    .X(_3198_));
 sky130_fd_sc_hd__nand2_1 _6610_ (.A(net203),
    .B(_3175_),
    .Y(_3199_));
 sky130_fd_sc_hd__o211a_1 _6611_ (.A1(_3196_),
    .A2(_3198_),
    .B1(_3199_),
    .C1(_3176_),
    .X(_3200_));
 sky130_fd_sc_hd__nor3_1 _6612_ (.A(_1157_),
    .B(_3194_),
    .C(_3200_),
    .Y(_0454_));
 sky130_fd_sc_hd__nor2_1 _6613_ (.A(\core_0.execute.alu_flag_reg.o_d[4] ),
    .B(_3176_),
    .Y(_3201_));
 sky130_fd_sc_hd__nand2_1 _6614_ (.A(_2582_),
    .B(_2611_),
    .Y(_3202_));
 sky130_fd_sc_hd__nand2_1 _6615_ (.A(_3177_),
    .B(_3202_),
    .Y(_3203_));
 sky130_fd_sc_hd__or2_1 _6616_ (.A(_2520_),
    .B(_2559_),
    .X(_3204_));
 sky130_fd_sc_hd__and2_1 _6617_ (.A(_3178_),
    .B(_3204_),
    .X(_3205_));
 sky130_fd_sc_hd__xor2_1 _6618_ (.A(_2338_),
    .B(_2364_),
    .X(_3206_));
 sky130_fd_sc_hd__xnor2_1 _6619_ (.A(_2456_),
    .B(_2491_),
    .Y(_3207_));
 sky130_fd_sc_hd__a21o_1 _6620_ (.A1(_2419_),
    .A2(_2424_),
    .B1(_2393_),
    .X(_3208_));
 sky130_fd_sc_hd__xnor2_1 _6621_ (.A(_2263_),
    .B(_2295_),
    .Y(_3209_));
 sky130_fd_sc_hd__xor2_1 _6622_ (.A(_2184_),
    .B(_2238_),
    .X(_3210_));
 sky130_fd_sc_hd__xnor2_1 _6623_ (.A(_1782_),
    .B(_2134_),
    .Y(_3211_));
 sky130_fd_sc_hd__xnor2_1 _6624_ (.A(_3210_),
    .B(_3211_),
    .Y(_3212_));
 sky130_fd_sc_hd__xnor2_1 _6625_ (.A(_3209_),
    .B(_3212_),
    .Y(_3213_));
 sky130_fd_sc_hd__a21o_1 _6626_ (.A1(_3179_),
    .A2(_3208_),
    .B1(_3213_),
    .X(_3214_));
 sky130_fd_sc_hd__nand3_1 _6627_ (.A(_3179_),
    .B(_3208_),
    .C(_3213_),
    .Y(_3215_));
 sky130_fd_sc_hd__nand3_1 _6628_ (.A(_3207_),
    .B(_3214_),
    .C(_3215_),
    .Y(_3216_));
 sky130_fd_sc_hd__a21o_1 _6629_ (.A1(_3214_),
    .A2(_3215_),
    .B1(_3207_),
    .X(_3217_));
 sky130_fd_sc_hd__nand3_1 _6630_ (.A(_3206_),
    .B(_3216_),
    .C(_3217_),
    .Y(_3218_));
 sky130_fd_sc_hd__a21o_1 _6631_ (.A1(_3216_),
    .A2(_3217_),
    .B1(_3206_),
    .X(_3219_));
 sky130_fd_sc_hd__nand3_1 _6632_ (.A(_3205_),
    .B(_3218_),
    .C(_3219_),
    .Y(_3220_));
 sky130_fd_sc_hd__a21o_1 _6633_ (.A1(_3218_),
    .A2(_3219_),
    .B1(_3205_),
    .X(_3221_));
 sky130_fd_sc_hd__and3_1 _6634_ (.A(_3203_),
    .B(_3220_),
    .C(_3221_),
    .X(_3222_));
 sky130_fd_sc_hd__a21oi_1 _6635_ (.A1(_3220_),
    .A2(_3221_),
    .B1(_3203_),
    .Y(_3223_));
 sky130_fd_sc_hd__nand2_1 _6636_ (.A(net204),
    .B(_3175_),
    .Y(_3224_));
 sky130_fd_sc_hd__o311a_1 _6637_ (.A1(_3175_),
    .A2(_3222_),
    .A3(_3223_),
    .B1(_3224_),
    .C1(_3176_),
    .X(_3225_));
 sky130_fd_sc_hd__nor3_1 _6638_ (.A(_1157_),
    .B(_3201_),
    .C(_3225_),
    .Y(_0455_));
 sky130_fd_sc_hd__mux2_1 _6639_ (.A0(net72),
    .A1(\core_0.execute.mem_stage_pc[0] ),
    .S(_1315_),
    .X(_3226_));
 sky130_fd_sc_hd__and2_1 _6640_ (.A(\core_0.dec_sreg_store ),
    .B(_2368_),
    .X(_3227_));
 sky130_fd_sc_hd__clkbuf_4 _6641_ (.A(_3227_),
    .X(_3228_));
 sky130_fd_sc_hd__buf_4 _6642_ (.A(_3228_),
    .X(_3229_));
 sky130_fd_sc_hd__mux2_1 _6643_ (.A0(_3226_),
    .A1(net194),
    .S(_3229_),
    .X(_3230_));
 sky130_fd_sc_hd__a21o_2 _6644_ (.A1(_1071_),
    .A2(_3228_),
    .B1(_0674_),
    .X(_3231_));
 sky130_fd_sc_hd__buf_4 _6645_ (.A(_3231_),
    .X(_3232_));
 sky130_fd_sc_hd__mux2_1 _6646_ (.A0(\core_0.execute.sreg_irq_pc.o_d[0] ),
    .A1(_3230_),
    .S(_3232_),
    .X(_3233_));
 sky130_fd_sc_hd__and2_1 _6647_ (.A(_1190_),
    .B(_3233_),
    .X(_3234_));
 sky130_fd_sc_hd__clkbuf_1 _6648_ (.A(_3234_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _6649_ (.A0(net79),
    .A1(\core_0.execute.mem_stage_pc[1] ),
    .S(_1315_),
    .X(_3235_));
 sky130_fd_sc_hd__mux2_1 _6650_ (.A0(_3235_),
    .A1(net201),
    .S(_3229_),
    .X(_3236_));
 sky130_fd_sc_hd__mux2_1 _6651_ (.A0(\core_0.execute.sreg_irq_pc.o_d[1] ),
    .A1(_3236_),
    .S(_3232_),
    .X(_3237_));
 sky130_fd_sc_hd__and2_1 _6652_ (.A(_1190_),
    .B(_3237_),
    .X(_3238_));
 sky130_fd_sc_hd__clkbuf_1 _6653_ (.A(_3238_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _6654_ (.A0(net80),
    .A1(\core_0.execute.mem_stage_pc[2] ),
    .S(_1315_),
    .X(_3239_));
 sky130_fd_sc_hd__mux2_1 _6655_ (.A0(_3239_),
    .A1(net202),
    .S(_3229_),
    .X(_3240_));
 sky130_fd_sc_hd__mux2_1 _6656_ (.A0(\core_0.execute.sreg_irq_pc.o_d[2] ),
    .A1(_3240_),
    .S(_3232_),
    .X(_3241_));
 sky130_fd_sc_hd__and2_1 _6657_ (.A(_1190_),
    .B(_3241_),
    .X(_3242_));
 sky130_fd_sc_hd__clkbuf_1 _6658_ (.A(_3242_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_4 _6659_ (.A(_0995_),
    .X(_3243_));
 sky130_fd_sc_hd__mux2_1 _6660_ (.A0(net81),
    .A1(\core_0.execute.mem_stage_pc[3] ),
    .S(_1315_),
    .X(_3244_));
 sky130_fd_sc_hd__mux2_1 _6661_ (.A0(_3244_),
    .A1(net203),
    .S(_3229_),
    .X(_3245_));
 sky130_fd_sc_hd__mux2_1 _6662_ (.A0(\core_0.execute.sreg_irq_pc.o_d[3] ),
    .A1(_3245_),
    .S(_3232_),
    .X(_3246_));
 sky130_fd_sc_hd__and2_1 _6663_ (.A(_3243_),
    .B(_3246_),
    .X(_3247_));
 sky130_fd_sc_hd__clkbuf_1 _6664_ (.A(_3247_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _6665_ (.A0(net82),
    .A1(\core_0.execute.mem_stage_pc[4] ),
    .S(_1315_),
    .X(_3248_));
 sky130_fd_sc_hd__mux2_1 _6666_ (.A0(_3248_),
    .A1(net204),
    .S(_3229_),
    .X(_3249_));
 sky130_fd_sc_hd__mux2_1 _6667_ (.A0(\core_0.execute.sreg_irq_pc.o_d[4] ),
    .A1(_3249_),
    .S(_3232_),
    .X(_3250_));
 sky130_fd_sc_hd__and2_1 _6668_ (.A(_3243_),
    .B(_3250_),
    .X(_3251_));
 sky130_fd_sc_hd__clkbuf_1 _6669_ (.A(_3251_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _6670_ (.A0(net83),
    .A1(\core_0.execute.mem_stage_pc[5] ),
    .S(_1315_),
    .X(_3252_));
 sky130_fd_sc_hd__mux2_1 _6671_ (.A0(_3252_),
    .A1(net205),
    .S(_3229_),
    .X(_3253_));
 sky130_fd_sc_hd__mux2_1 _6672_ (.A0(\core_0.execute.sreg_irq_pc.o_d[5] ),
    .A1(_3253_),
    .S(_3232_),
    .X(_3254_));
 sky130_fd_sc_hd__and2_1 _6673_ (.A(_3243_),
    .B(_3254_),
    .X(_3255_));
 sky130_fd_sc_hd__clkbuf_1 _6674_ (.A(_3255_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _6675_ (.A0(net84),
    .A1(\core_0.execute.mem_stage_pc[6] ),
    .S(_1315_),
    .X(_3256_));
 sky130_fd_sc_hd__mux2_1 _6676_ (.A0(_3256_),
    .A1(net206),
    .S(_3229_),
    .X(_3257_));
 sky130_fd_sc_hd__mux2_1 _6677_ (.A0(\core_0.execute.sreg_irq_pc.o_d[6] ),
    .A1(_3257_),
    .S(_3232_),
    .X(_3258_));
 sky130_fd_sc_hd__and2_1 _6678_ (.A(_3243_),
    .B(_3258_),
    .X(_3259_));
 sky130_fd_sc_hd__clkbuf_1 _6679_ (.A(_3259_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _6680_ (.A0(net85),
    .A1(\core_0.execute.mem_stage_pc[7] ),
    .S(_1315_),
    .X(_3260_));
 sky130_fd_sc_hd__mux2_1 _6681_ (.A0(_3260_),
    .A1(net207),
    .S(_3229_),
    .X(_3261_));
 sky130_fd_sc_hd__mux2_1 _6682_ (.A0(\core_0.execute.sreg_irq_pc.o_d[7] ),
    .A1(_3261_),
    .S(_3232_),
    .X(_3262_));
 sky130_fd_sc_hd__and2_1 _6683_ (.A(_3243_),
    .B(_3262_),
    .X(_3263_));
 sky130_fd_sc_hd__clkbuf_1 _6684_ (.A(_3263_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _6685_ (.A0(net86),
    .A1(\core_0.execute.mem_stage_pc[8] ),
    .S(net37),
    .X(_3264_));
 sky130_fd_sc_hd__mux2_1 _6686_ (.A0(_3264_),
    .A1(net208),
    .S(_3229_),
    .X(_3265_));
 sky130_fd_sc_hd__mux2_1 _6687_ (.A0(\core_0.execute.sreg_irq_pc.o_d[8] ),
    .A1(_3265_),
    .S(_3232_),
    .X(_3266_));
 sky130_fd_sc_hd__and2_1 _6688_ (.A(_3243_),
    .B(_3266_),
    .X(_3267_));
 sky130_fd_sc_hd__clkbuf_1 _6689_ (.A(_3267_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _6690_ (.A0(net87),
    .A1(\core_0.execute.mem_stage_pc[9] ),
    .S(net37),
    .X(_3268_));
 sky130_fd_sc_hd__mux2_1 _6691_ (.A0(_3268_),
    .A1(net209),
    .S(_3229_),
    .X(_3269_));
 sky130_fd_sc_hd__mux2_1 _6692_ (.A0(\core_0.execute.sreg_irq_pc.o_d[9] ),
    .A1(_3269_),
    .S(_3232_),
    .X(_3270_));
 sky130_fd_sc_hd__and2_1 _6693_ (.A(_3243_),
    .B(_3270_),
    .X(_3271_));
 sky130_fd_sc_hd__clkbuf_1 _6694_ (.A(_3271_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _6695_ (.A0(net73),
    .A1(\core_0.execute.mem_stage_pc[10] ),
    .S(net37),
    .X(_3272_));
 sky130_fd_sc_hd__mux2_1 _6696_ (.A0(_3272_),
    .A1(net195),
    .S(_3228_),
    .X(_3273_));
 sky130_fd_sc_hd__mux2_1 _6697_ (.A0(\core_0.execute.sreg_irq_pc.o_d[10] ),
    .A1(_3273_),
    .S(_3231_),
    .X(_3274_));
 sky130_fd_sc_hd__and2_1 _6698_ (.A(_3243_),
    .B(_3274_),
    .X(_3275_));
 sky130_fd_sc_hd__clkbuf_1 _6699_ (.A(_3275_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _6700_ (.A0(net74),
    .A1(\core_0.execute.mem_stage_pc[11] ),
    .S(net37),
    .X(_3276_));
 sky130_fd_sc_hd__mux2_1 _6701_ (.A0(_3276_),
    .A1(net196),
    .S(_3228_),
    .X(_3277_));
 sky130_fd_sc_hd__mux2_1 _6702_ (.A0(\core_0.execute.sreg_irq_pc.o_d[11] ),
    .A1(_3277_),
    .S(_3231_),
    .X(_3278_));
 sky130_fd_sc_hd__and2_1 _6703_ (.A(_3243_),
    .B(_3278_),
    .X(_3279_));
 sky130_fd_sc_hd__clkbuf_1 _6704_ (.A(_3279_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _6705_ (.A0(net75),
    .A1(\core_0.execute.mem_stage_pc[12] ),
    .S(net37),
    .X(_3280_));
 sky130_fd_sc_hd__mux2_1 _6706_ (.A0(_3280_),
    .A1(net197),
    .S(_3228_),
    .X(_3281_));
 sky130_fd_sc_hd__mux2_1 _6707_ (.A0(\core_0.execute.sreg_irq_pc.o_d[12] ),
    .A1(_3281_),
    .S(_3231_),
    .X(_3282_));
 sky130_fd_sc_hd__and2_1 _6708_ (.A(_3243_),
    .B(_3282_),
    .X(_3283_));
 sky130_fd_sc_hd__clkbuf_1 _6709_ (.A(_3283_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_4 _6710_ (.A(_0995_),
    .X(_3284_));
 sky130_fd_sc_hd__mux2_1 _6711_ (.A0(net76),
    .A1(\core_0.execute.mem_stage_pc[13] ),
    .S(net37),
    .X(_3285_));
 sky130_fd_sc_hd__mux2_1 _6712_ (.A0(_3285_),
    .A1(net198),
    .S(_3228_),
    .X(_3286_));
 sky130_fd_sc_hd__mux2_1 _6713_ (.A0(\core_0.execute.sreg_irq_pc.o_d[13] ),
    .A1(_3286_),
    .S(_3231_),
    .X(_3287_));
 sky130_fd_sc_hd__and2_1 _6714_ (.A(_3284_),
    .B(_3287_),
    .X(_3288_));
 sky130_fd_sc_hd__clkbuf_1 _6715_ (.A(_3288_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _6716_ (.A0(net77),
    .A1(\core_0.execute.mem_stage_pc[14] ),
    .S(net37),
    .X(_3289_));
 sky130_fd_sc_hd__mux2_1 _6717_ (.A0(_3289_),
    .A1(net199),
    .S(_3228_),
    .X(_3290_));
 sky130_fd_sc_hd__mux2_1 _6718_ (.A0(\core_0.execute.sreg_irq_pc.o_d[14] ),
    .A1(_3290_),
    .S(_3231_),
    .X(_3291_));
 sky130_fd_sc_hd__and2_1 _6719_ (.A(_3284_),
    .B(_3291_),
    .X(_3292_));
 sky130_fd_sc_hd__clkbuf_1 _6720_ (.A(_3292_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _6721_ (.A0(net78),
    .A1(\core_0.execute.mem_stage_pc[15] ),
    .S(net37),
    .X(_3293_));
 sky130_fd_sc_hd__mux2_1 _6722_ (.A0(_3293_),
    .A1(net200),
    .S(_3228_),
    .X(_3294_));
 sky130_fd_sc_hd__mux2_1 _6723_ (.A0(\core_0.execute.sreg_irq_pc.o_d[15] ),
    .A1(_3294_),
    .S(_3231_),
    .X(_3295_));
 sky130_fd_sc_hd__and2_1 _6724_ (.A(_3284_),
    .B(_3295_),
    .X(_3296_));
 sky130_fd_sc_hd__clkbuf_1 _6725_ (.A(_3296_),
    .X(_0471_));
 sky130_fd_sc_hd__and3_1 _6726_ (.A(\core_0.execute.sreg_priv_control.o_d[0] ),
    .B(_1152_),
    .C(_0746_),
    .X(_3297_));
 sky130_fd_sc_hd__and3_1 _6727_ (.A(_3297_),
    .B(_2064_),
    .C(_2066_),
    .X(_3298_));
 sky130_fd_sc_hd__nor2_1 _6728_ (.A(_0674_),
    .B(_3298_),
    .Y(_3299_));
 sky130_fd_sc_hd__a221o_1 _6729_ (.A1(net194),
    .A2(_3298_),
    .B1(_3299_),
    .B2(\core_0.execute.sreg_jtr_buff.o_d[0] ),
    .C1(_1157_),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _6730_ (.A1(net201),
    .A2(_3298_),
    .B1(_3299_),
    .B2(\core_0.execute.sreg_jtr_buff.o_d[1] ),
    .X(_3300_));
 sky130_fd_sc_hd__and2_1 _6731_ (.A(_3284_),
    .B(_3300_),
    .X(_3301_));
 sky130_fd_sc_hd__clkbuf_1 _6732_ (.A(_3301_),
    .X(_0473_));
 sky130_fd_sc_hd__a22o_1 _6733_ (.A1(net202),
    .A2(_3298_),
    .B1(_3299_),
    .B2(\core_0.execute.sreg_jtr_buff.o_d[2] ),
    .X(_3302_));
 sky130_fd_sc_hd__and2_1 _6734_ (.A(_3284_),
    .B(_3302_),
    .X(_3303_));
 sky130_fd_sc_hd__clkbuf_1 _6735_ (.A(_3303_),
    .X(_0474_));
 sky130_fd_sc_hd__nor2_1 _6736_ (.A(_0674_),
    .B(_1040_),
    .Y(_3304_));
 sky130_fd_sc_hd__a221o_1 _6737_ (.A1(\core_0.execute.sreg_jtr_buff.o_d[0] ),
    .A2(_1040_),
    .B1(_3304_),
    .B2(net106),
    .C1(_1157_),
    .X(_0475_));
 sky130_fd_sc_hd__a22o_1 _6738_ (.A1(\core_0.execute.sreg_jtr_buff.o_d[1] ),
    .A2(_1040_),
    .B1(_3304_),
    .B2(\core_0.execute.trap_flag ),
    .X(_3305_));
 sky130_fd_sc_hd__and2_1 _6739_ (.A(_3284_),
    .B(_3305_),
    .X(_3306_));
 sky130_fd_sc_hd__clkbuf_1 _6740_ (.A(_3306_),
    .X(_0476_));
 sky130_fd_sc_hd__a22o_1 _6741_ (.A1(\core_0.execute.sreg_jtr_buff.o_d[2] ),
    .A2(_1040_),
    .B1(_3304_),
    .B2(_0675_),
    .X(_3307_));
 sky130_fd_sc_hd__and2_1 _6742_ (.A(_3284_),
    .B(_3307_),
    .X(_3308_));
 sky130_fd_sc_hd__clkbuf_1 _6743_ (.A(_3308_),
    .X(_0477_));
 sky130_fd_sc_hd__and3_1 _6744_ (.A(_1152_),
    .B(_1071_),
    .C(_2369_),
    .X(_3309_));
 sky130_fd_sc_hd__clkbuf_4 _6745_ (.A(_3309_),
    .X(_3310_));
 sky130_fd_sc_hd__clkbuf_4 _6746_ (.A(_3310_),
    .X(_3311_));
 sky130_fd_sc_hd__clkbuf_4 _6747_ (.A(_3309_),
    .X(_3312_));
 sky130_fd_sc_hd__nand2_1 _6748_ (.A(_0664_),
    .B(_3312_),
    .Y(_3313_));
 sky130_fd_sc_hd__o211a_1 _6749_ (.A1(\core_0.execute.sreg_scratch.o_d[0] ),
    .A2(_3311_),
    .B1(_3313_),
    .C1(_2861_),
    .X(_0478_));
 sky130_fd_sc_hd__a21oi_1 _6750_ (.A1(_0655_),
    .A2(_3310_),
    .B1(_1157_),
    .Y(_3314_));
 sky130_fd_sc_hd__o21a_1 _6751_ (.A1(\core_0.execute.sreg_scratch.o_d[1] ),
    .A2(_3311_),
    .B1(_3314_),
    .X(_0479_));
 sky130_fd_sc_hd__inv_2 _6752_ (.A(net202),
    .Y(_3315_));
 sky130_fd_sc_hd__o21ai_1 _6753_ (.A1(\core_0.execute.sreg_scratch.o_d[2] ),
    .A2(_3310_),
    .B1(_1075_),
    .Y(_3316_));
 sky130_fd_sc_hd__a21oi_1 _6754_ (.A1(_3315_),
    .A2(_3312_),
    .B1(_3316_),
    .Y(_0480_));
 sky130_fd_sc_hd__nand2_1 _6755_ (.A(_0639_),
    .B(_3312_),
    .Y(_3317_));
 sky130_fd_sc_hd__clkbuf_4 _6756_ (.A(_0996_),
    .X(_3318_));
 sky130_fd_sc_hd__o211a_1 _6757_ (.A1(\core_0.execute.sreg_scratch.o_d[3] ),
    .A2(_3311_),
    .B1(_3317_),
    .C1(_3318_),
    .X(_0481_));
 sky130_fd_sc_hd__nand2_1 _6758_ (.A(_0633_),
    .B(_3312_),
    .Y(_3319_));
 sky130_fd_sc_hd__o211a_1 _6759_ (.A1(\core_0.execute.sreg_scratch.o_d[4] ),
    .A2(_3311_),
    .B1(_3319_),
    .C1(_3318_),
    .X(_0482_));
 sky130_fd_sc_hd__nand2_1 _6760_ (.A(_0627_),
    .B(_3312_),
    .Y(_3320_));
 sky130_fd_sc_hd__o211a_1 _6761_ (.A1(\core_0.execute.sreg_scratch.o_d[5] ),
    .A2(_3311_),
    .B1(_3320_),
    .C1(_3318_),
    .X(_0483_));
 sky130_fd_sc_hd__inv_2 _6762_ (.A(net206),
    .Y(_3321_));
 sky130_fd_sc_hd__o21ai_1 _6763_ (.A1(\core_0.execute.sreg_scratch.o_d[6] ),
    .A2(_3310_),
    .B1(_1075_),
    .Y(_3322_));
 sky130_fd_sc_hd__a21oi_1 _6764_ (.A1(_3321_),
    .A2(_3312_),
    .B1(_3322_),
    .Y(_0484_));
 sky130_fd_sc_hd__nand2_1 _6765_ (.A(_0613_),
    .B(_3310_),
    .Y(_3323_));
 sky130_fd_sc_hd__o211a_1 _6766_ (.A1(\core_0.execute.sreg_scratch.o_d[7] ),
    .A2(_3311_),
    .B1(_3323_),
    .C1(_3318_),
    .X(_0485_));
 sky130_fd_sc_hd__nand2_1 _6767_ (.A(_0604_),
    .B(_3310_),
    .Y(_3324_));
 sky130_fd_sc_hd__o211a_1 _6768_ (.A1(\core_0.execute.sreg_scratch.o_d[8] ),
    .A2(_3311_),
    .B1(_3324_),
    .C1(_3318_),
    .X(_0486_));
 sky130_fd_sc_hd__nand2_1 _6769_ (.A(_0598_),
    .B(_3310_),
    .Y(_3325_));
 sky130_fd_sc_hd__o211a_1 _6770_ (.A1(\core_0.execute.sreg_scratch.o_d[9] ),
    .A2(_3311_),
    .B1(_3325_),
    .C1(_3318_),
    .X(_0487_));
 sky130_fd_sc_hd__nand2_1 _6771_ (.A(_0592_),
    .B(_3310_),
    .Y(_3326_));
 sky130_fd_sc_hd__o211a_1 _6772_ (.A1(\core_0.execute.sreg_scratch.o_d[10] ),
    .A2(_3311_),
    .B1(_3326_),
    .C1(_3318_),
    .X(_0488_));
 sky130_fd_sc_hd__o21ai_1 _6773_ (.A1(\core_0.execute.sreg_scratch.o_d[11] ),
    .A2(_3310_),
    .B1(_1075_),
    .Y(_3327_));
 sky130_fd_sc_hd__a21oi_1 _6774_ (.A1(_1340_),
    .A2(_3312_),
    .B1(_3327_),
    .Y(_0489_));
 sky130_fd_sc_hd__nand2_1 _6775_ (.A(_0579_),
    .B(_3310_),
    .Y(_3328_));
 sky130_fd_sc_hd__o211a_1 _6776_ (.A1(\core_0.execute.sreg_scratch.o_d[12] ),
    .A2(_3311_),
    .B1(_3328_),
    .C1(_3318_),
    .X(_0490_));
 sky130_fd_sc_hd__or2b_1 _6777_ (.A(net198),
    .B_N(_3309_),
    .X(_3329_));
 sky130_fd_sc_hd__o211a_1 _6778_ (.A1(\core_0.execute.sreg_scratch.o_d[13] ),
    .A2(_3312_),
    .B1(_3329_),
    .C1(_3318_),
    .X(_0491_));
 sky130_fd_sc_hd__or2b_1 _6779_ (.A(net199),
    .B_N(_3309_),
    .X(_3330_));
 sky130_fd_sc_hd__o211a_1 _6780_ (.A1(\core_0.execute.sreg_scratch.o_d[14] ),
    .A2(_3312_),
    .B1(_3330_),
    .C1(_3318_),
    .X(_0492_));
 sky130_fd_sc_hd__or2b_1 _6781_ (.A(net200),
    .B_N(_3309_),
    .X(_3331_));
 sky130_fd_sc_hd__clkbuf_4 _6782_ (.A(_0996_),
    .X(_3332_));
 sky130_fd_sc_hd__o211a_1 _6783_ (.A1(\core_0.execute.sreg_scratch.o_d[15] ),
    .A2(_3312_),
    .B1(_3331_),
    .C1(_3332_),
    .X(_0493_));
 sky130_fd_sc_hd__a32o_1 _6784_ (.A1(\core_0.execute.irq_en ),
    .A2(net18),
    .A3(_1075_),
    .B1(_2870_),
    .B2(\core_0.execute.sreg_irq_flags.o_d[0] ),
    .X(_0494_));
 sky130_fd_sc_hd__inv_2 _6785_ (.A(\core_0.execute.sreg_irq_flags.o_d[1] ),
    .Y(_3333_));
 sky130_fd_sc_hd__nor2_1 _6786_ (.A(_3333_),
    .B(_0672_),
    .Y(_3334_));
 sky130_fd_sc_hd__o21a_1 _6787_ (.A1(\core_0.execute.prev_sys ),
    .A2(_3334_),
    .B1(_0997_),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_1 _6788_ (.A1(\core_0.execute.sreg_irq_flags.i_d[2] ),
    .A2(_1075_),
    .B1(_2870_),
    .B2(\core_0.execute.sreg_irq_flags.o_d[2] ),
    .X(_0496_));
 sky130_fd_sc_hd__a22o_1 _6789_ (.A1(_1315_),
    .A2(_1075_),
    .B1(_2870_),
    .B2(\core_0.execute.sreg_irq_flags.o_d[3] ),
    .X(_0497_));
 sky130_fd_sc_hd__a32o_1 _6790_ (.A1(\core_0.execute.irq_en ),
    .A2(net19),
    .A3(_1075_),
    .B1(_2870_),
    .B2(\core_0.execute.sreg_irq_flags.o_d[4] ),
    .X(_0498_));
 sky130_fd_sc_hd__and2_1 _6791_ (.A(\core_0.dec_sreg_store ),
    .B(_2075_),
    .X(_3335_));
 sky130_fd_sc_hd__and2_2 _6792_ (.A(_0675_),
    .B(_1040_),
    .X(_3336_));
 sky130_fd_sc_hd__and3_1 _6793_ (.A(_0675_),
    .B(net77),
    .C(_1687_),
    .X(_3337_));
 sky130_fd_sc_hd__o31a_1 _6794_ (.A1(_3335_),
    .A2(_3336_),
    .A3(_3337_),
    .B1(_0746_),
    .X(_3338_));
 sky130_fd_sc_hd__clkbuf_4 _6795_ (.A(_3338_),
    .X(_3339_));
 sky130_fd_sc_hd__nor2_1 _6796_ (.A(\core_0.execute.pc_high_out[0] ),
    .B(_3339_),
    .Y(_3340_));
 sky130_fd_sc_hd__nand2_4 _6797_ (.A(_1152_),
    .B(_2075_),
    .Y(_3341_));
 sky130_fd_sc_hd__nand2_4 _6798_ (.A(_0675_),
    .B(_1040_),
    .Y(_3342_));
 sky130_fd_sc_hd__nor2_1 _6799_ (.A(\core_0.execute.pc_high_buff_out[0] ),
    .B(_3342_),
    .Y(_3343_));
 sky130_fd_sc_hd__a211o_1 _6800_ (.A1(\core_0.execute.pc_high_out[0] ),
    .A2(_3342_),
    .B1(_3343_),
    .C1(_3335_),
    .X(_3344_));
 sky130_fd_sc_hd__o211a_1 _6801_ (.A1(_0664_),
    .A2(_3341_),
    .B1(_3339_),
    .C1(_3344_),
    .X(_3345_));
 sky130_fd_sc_hd__nor3_1 _6802_ (.A(_1157_),
    .B(_3340_),
    .C(_3345_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _6803_ (.A(\core_0.execute.pc_high_out[1] ),
    .B(\core_0.execute.pc_high_out[0] ),
    .Y(_3346_));
 sky130_fd_sc_hd__o21a_1 _6804_ (.A1(\core_0.execute.pc_high_out[1] ),
    .A2(\core_0.execute.pc_high_out[0] ),
    .B1(_3342_),
    .X(_3347_));
 sky130_fd_sc_hd__a22o_1 _6805_ (.A1(\core_0.execute.pc_high_buff_out[1] ),
    .A2(_3336_),
    .B1(_3346_),
    .B2(_3347_),
    .X(_3348_));
 sky130_fd_sc_hd__mux2_1 _6806_ (.A0(net201),
    .A1(_3348_),
    .S(_3341_),
    .X(_3349_));
 sky130_fd_sc_hd__mux2_1 _6807_ (.A0(\core_0.execute.pc_high_out[1] ),
    .A1(_3349_),
    .S(_3339_),
    .X(_3350_));
 sky130_fd_sc_hd__and2_1 _6808_ (.A(_3284_),
    .B(_3350_),
    .X(_3351_));
 sky130_fd_sc_hd__clkbuf_1 _6809_ (.A(_3351_),
    .X(_0500_));
 sky130_fd_sc_hd__xnor2_1 _6810_ (.A(\core_0.execute.pc_high_out[2] ),
    .B(_3346_),
    .Y(_3352_));
 sky130_fd_sc_hd__mux2_1 _6811_ (.A0(\core_0.execute.pc_high_buff_out[2] ),
    .A1(_3352_),
    .S(_3342_),
    .X(_3353_));
 sky130_fd_sc_hd__mux2_1 _6812_ (.A0(net202),
    .A1(_3353_),
    .S(_3341_),
    .X(_3354_));
 sky130_fd_sc_hd__mux2_1 _6813_ (.A0(\core_0.execute.pc_high_out[2] ),
    .A1(_3354_),
    .S(_3339_),
    .X(_3355_));
 sky130_fd_sc_hd__and2_1 _6814_ (.A(_3284_),
    .B(_3355_),
    .X(_3356_));
 sky130_fd_sc_hd__clkbuf_1 _6815_ (.A(_3356_),
    .X(_0501_));
 sky130_fd_sc_hd__and4_1 _6816_ (.A(\core_0.execute.pc_high_out[3] ),
    .B(\core_0.execute.pc_high_out[2] ),
    .C(\core_0.execute.pc_high_out[1] ),
    .D(\core_0.execute.pc_high_out[0] ),
    .X(_3357_));
 sky130_fd_sc_hd__a31o_1 _6817_ (.A1(\core_0.execute.pc_high_out[2] ),
    .A2(\core_0.execute.pc_high_out[1] ),
    .A3(\core_0.execute.pc_high_out[0] ),
    .B1(\core_0.execute.pc_high_out[3] ),
    .X(_3358_));
 sky130_fd_sc_hd__nand2_1 _6818_ (.A(_3342_),
    .B(_3358_),
    .Y(_3359_));
 sky130_fd_sc_hd__a2bb2o_1 _6819_ (.A1_N(_3357_),
    .A2_N(_3359_),
    .B1(\core_0.execute.pc_high_buff_out[3] ),
    .B2(_3336_),
    .X(_3360_));
 sky130_fd_sc_hd__mux2_1 _6820_ (.A0(net203),
    .A1(_3360_),
    .S(_3341_),
    .X(_3361_));
 sky130_fd_sc_hd__mux2_1 _6821_ (.A0(\core_0.execute.pc_high_out[3] ),
    .A1(_3361_),
    .S(_3339_),
    .X(_3362_));
 sky130_fd_sc_hd__and2_1 _6822_ (.A(_3284_),
    .B(_3362_),
    .X(_3363_));
 sky130_fd_sc_hd__clkbuf_1 _6823_ (.A(_3363_),
    .X(_0502_));
 sky130_fd_sc_hd__o21ai_1 _6824_ (.A1(\core_0.execute.pc_high_out[4] ),
    .A2(_3357_),
    .B1(_3342_),
    .Y(_3364_));
 sky130_fd_sc_hd__a21oi_1 _6825_ (.A1(\core_0.execute.pc_high_out[4] ),
    .A2(_3357_),
    .B1(_3364_),
    .Y(_3365_));
 sky130_fd_sc_hd__a21oi_1 _6826_ (.A1(\core_0.execute.pc_high_buff_out[4] ),
    .A2(_3336_),
    .B1(_3365_),
    .Y(_3366_));
 sky130_fd_sc_hd__mux2_1 _6827_ (.A0(_0633_),
    .A1(_3366_),
    .S(_3341_),
    .X(_3367_));
 sky130_fd_sc_hd__nand2_1 _6828_ (.A(_3339_),
    .B(_3367_),
    .Y(_3368_));
 sky130_fd_sc_hd__o211a_1 _6829_ (.A1(\core_0.execute.pc_high_out[4] ),
    .A2(_3339_),
    .B1(_3368_),
    .C1(_3332_),
    .X(_0503_));
 sky130_fd_sc_hd__and3_1 _6830_ (.A(\core_0.execute.pc_high_out[5] ),
    .B(\core_0.execute.pc_high_out[4] ),
    .C(_3357_),
    .X(_3369_));
 sky130_fd_sc_hd__a21oi_1 _6831_ (.A1(\core_0.execute.pc_high_out[4] ),
    .A2(_3357_),
    .B1(\core_0.execute.pc_high_out[5] ),
    .Y(_3370_));
 sky130_fd_sc_hd__o21ai_1 _6832_ (.A1(_3369_),
    .A2(_3370_),
    .B1(_3342_),
    .Y(_3371_));
 sky130_fd_sc_hd__o211ai_1 _6833_ (.A1(\core_0.execute.pc_high_buff_out[5] ),
    .A2(_3342_),
    .B1(_3371_),
    .C1(_3341_),
    .Y(_3372_));
 sky130_fd_sc_hd__o211ai_1 _6834_ (.A1(_0627_),
    .A2(_3341_),
    .B1(_3339_),
    .C1(_3372_),
    .Y(_3373_));
 sky130_fd_sc_hd__o211a_1 _6835_ (.A1(\core_0.execute.pc_high_out[5] ),
    .A2(_3339_),
    .B1(_3373_),
    .C1(_3332_),
    .X(_0504_));
 sky130_fd_sc_hd__nand2_1 _6836_ (.A(\core_0.execute.pc_high_out[6] ),
    .B(_3369_),
    .Y(_3374_));
 sky130_fd_sc_hd__o21a_1 _6837_ (.A1(\core_0.execute.pc_high_out[6] ),
    .A2(_3369_),
    .B1(_3342_),
    .X(_3375_));
 sky130_fd_sc_hd__a22o_1 _6838_ (.A1(\core_0.execute.pc_high_buff_out[6] ),
    .A2(_3336_),
    .B1(_3374_),
    .B2(_3375_),
    .X(_3376_));
 sky130_fd_sc_hd__mux2_1 _6839_ (.A0(net206),
    .A1(_3376_),
    .S(_3341_),
    .X(_3377_));
 sky130_fd_sc_hd__mux2_1 _6840_ (.A0(\core_0.execute.pc_high_out[6] ),
    .A1(_3377_),
    .S(_3339_),
    .X(_3378_));
 sky130_fd_sc_hd__and2_1 _6841_ (.A(_1314_),
    .B(_3378_),
    .X(_3379_));
 sky130_fd_sc_hd__clkbuf_1 _6842_ (.A(_3379_),
    .X(_0505_));
 sky130_fd_sc_hd__xnor2_1 _6843_ (.A(\core_0.execute.pc_high_out[7] ),
    .B(_3374_),
    .Y(_3380_));
 sky130_fd_sc_hd__mux2_1 _6844_ (.A0(\core_0.execute.pc_high_buff_out[7] ),
    .A1(_3380_),
    .S(_3342_),
    .X(_3381_));
 sky130_fd_sc_hd__mux2_1 _6845_ (.A0(net207),
    .A1(_3381_),
    .S(_3341_),
    .X(_3382_));
 sky130_fd_sc_hd__mux2_1 _6846_ (.A0(\core_0.execute.pc_high_out[7] ),
    .A1(_3382_),
    .S(_3338_),
    .X(_3383_));
 sky130_fd_sc_hd__or2_1 _6847_ (.A(_1122_),
    .B(_3383_),
    .X(_3384_));
 sky130_fd_sc_hd__clkbuf_1 _6848_ (.A(_3384_),
    .X(_0506_));
 sky130_fd_sc_hd__a22o_1 _6849_ (.A1(_0675_),
    .A2(\core_0.dec_sreg_jal_over ),
    .B1(_1152_),
    .B2(_2072_),
    .X(_3385_));
 sky130_fd_sc_hd__and2_1 _6850_ (.A(_0746_),
    .B(_3385_),
    .X(_3386_));
 sky130_fd_sc_hd__clkbuf_2 _6851_ (.A(_3386_),
    .X(_3387_));
 sky130_fd_sc_hd__buf_2 _6852_ (.A(_3387_),
    .X(_3388_));
 sky130_fd_sc_hd__and4_1 _6853_ (.A(net178),
    .B(_1033_),
    .C(_1034_),
    .D(_2071_),
    .X(_3389_));
 sky130_fd_sc_hd__nand2_4 _6854_ (.A(_1152_),
    .B(_3389_),
    .Y(_3390_));
 sky130_fd_sc_hd__mux2_1 _6855_ (.A0(_0664_),
    .A1(_0689_),
    .S(_3390_),
    .X(_3391_));
 sky130_fd_sc_hd__nand2_1 _6856_ (.A(_3388_),
    .B(_3391_),
    .Y(_3392_));
 sky130_fd_sc_hd__o211a_1 _6857_ (.A1(\core_0.execute.pc_high_buff_out[0] ),
    .A2(_3388_),
    .B1(_3392_),
    .C1(_3332_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _6858_ (.A0(_0655_),
    .A1(_0687_),
    .S(_3390_),
    .X(_3393_));
 sky130_fd_sc_hd__nand2_1 _6859_ (.A(_3388_),
    .B(_3393_),
    .Y(_3394_));
 sky130_fd_sc_hd__o211a_1 _6860_ (.A1(\core_0.execute.pc_high_buff_out[1] ),
    .A2(_3388_),
    .B1(_3394_),
    .C1(_3332_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _6861_ (.A0(_3315_),
    .A1(_0676_),
    .S(_3390_),
    .X(_3395_));
 sky130_fd_sc_hd__nand2_1 _6862_ (.A(_3388_),
    .B(_3395_),
    .Y(_3396_));
 sky130_fd_sc_hd__o211a_1 _6863_ (.A1(\core_0.execute.pc_high_buff_out[2] ),
    .A2(_3388_),
    .B1(_3396_),
    .C1(_3332_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _6864_ (.A0(_0639_),
    .A1(_0678_),
    .S(_3390_),
    .X(_3397_));
 sky130_fd_sc_hd__nand2_1 _6865_ (.A(_3387_),
    .B(_3397_),
    .Y(_3398_));
 sky130_fd_sc_hd__o211a_1 _6866_ (.A1(\core_0.execute.pc_high_buff_out[3] ),
    .A2(_3388_),
    .B1(_3398_),
    .C1(_3332_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _6867_ (.A0(_0633_),
    .A1(_0682_),
    .S(_3390_),
    .X(_3399_));
 sky130_fd_sc_hd__nand2_1 _6868_ (.A(_3387_),
    .B(_3399_),
    .Y(_3400_));
 sky130_fd_sc_hd__o211a_1 _6869_ (.A1(\core_0.execute.pc_high_buff_out[4] ),
    .A2(_3388_),
    .B1(_3400_),
    .C1(_3332_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _6870_ (.A0(_0627_),
    .A1(_0685_),
    .S(_3390_),
    .X(_3401_));
 sky130_fd_sc_hd__nand2_1 _6871_ (.A(_3387_),
    .B(_3401_),
    .Y(_3402_));
 sky130_fd_sc_hd__o211a_1 _6872_ (.A1(\core_0.execute.pc_high_buff_out[5] ),
    .A2(_3388_),
    .B1(_3402_),
    .C1(_3332_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _6873_ (.A0(_3321_),
    .A1(_0681_),
    .S(_3390_),
    .X(_3403_));
 sky130_fd_sc_hd__nand2_1 _6874_ (.A(_3387_),
    .B(_3403_),
    .Y(_3404_));
 sky130_fd_sc_hd__o211a_1 _6875_ (.A1(\core_0.execute.pc_high_buff_out[6] ),
    .A2(_3388_),
    .B1(_3404_),
    .C1(_3332_),
    .X(_0513_));
 sky130_fd_sc_hd__clkinv_2 _6876_ (.A(\core_0.execute.pc_high_buff_out[7] ),
    .Y(_3405_));
 sky130_fd_sc_hd__mux2_1 _6877_ (.A0(_0613_),
    .A1(_0677_),
    .S(_3390_),
    .X(_3406_));
 sky130_fd_sc_hd__mux2_1 _6878_ (.A0(_3405_),
    .A1(_3406_),
    .S(_3387_),
    .X(_3407_));
 sky130_fd_sc_hd__nand2_1 _6879_ (.A(_0997_),
    .B(_3407_),
    .Y(_0514_));
 sky130_fd_sc_hd__dfxtp_4 _6880_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0015_),
    .Q(\core_0.decode.o_submit ));
 sky130_fd_sc_hd__dfxtp_2 _6881_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0016_),
    .Q(\core_0.dec_pc_inc ));
 sky130_fd_sc_hd__dfxtp_2 _6882_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0017_),
    .Q(\core_0.dec_r_bus_imm ));
 sky130_fd_sc_hd__dfxtp_1 _6883_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0018_),
    .Q(\core_0.dec_alu_flags_ie ));
 sky130_fd_sc_hd__dfxtp_1 _6884_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0019_),
    .Q(\core_0.dec_alu_carry_en ));
 sky130_fd_sc_hd__dfxtp_1 _6885_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0020_),
    .Q(\core_0.dec_l_reg_sel[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6886_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0021_),
    .Q(\core_0.dec_l_reg_sel[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6887_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0022_),
    .Q(\core_0.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6888_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0023_),
    .Q(\core_0.dec_r_reg_sel[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6889_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0024_),
    .Q(\core_0.dec_r_reg_sel[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6890_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0025_),
    .Q(\core_0.dec_r_reg_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6891_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0026_),
    .Q(\core_0.dec_rf_ie[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6892_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0027_),
    .Q(\core_0.dec_rf_ie[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6893_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0028_),
    .Q(\core_0.dec_rf_ie[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6894_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0029_),
    .Q(\core_0.dec_rf_ie[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6895_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0030_),
    .Q(\core_0.dec_rf_ie[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6896_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0031_),
    .Q(\core_0.dec_rf_ie[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6897_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0032_),
    .Q(\core_0.dec_rf_ie[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6898_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0033_),
    .Q(\core_0.dec_rf_ie[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6899_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0034_),
    .Q(\core_0.dec_jump_cond_code[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6900_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0035_),
    .Q(\core_0.dec_jump_cond_code[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6901_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0036_),
    .Q(\core_0.dec_jump_cond_code[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6902_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0037_),
    .Q(\core_0.dec_jump_cond_code[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6903_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0038_),
    .Q(\core_0.dec_jump_cond_code[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6904_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0039_),
    .Q(net178));
 sky130_fd_sc_hd__dfxtp_4 _6905_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0040_),
    .Q(net185));
 sky130_fd_sc_hd__dfxtp_4 _6906_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0041_),
    .Q(net186));
 sky130_fd_sc_hd__dfxtp_4 _6907_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0042_),
    .Q(net187));
 sky130_fd_sc_hd__dfxtp_4 _6908_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0043_),
    .Q(net188));
 sky130_fd_sc_hd__dfxtp_4 _6909_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0044_),
    .Q(net189));
 sky130_fd_sc_hd__dfxtp_4 _6910_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0045_),
    .Q(net190));
 sky130_fd_sc_hd__dfxtp_4 _6911_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0046_),
    .Q(net191));
 sky130_fd_sc_hd__dfxtp_4 _6912_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0047_),
    .Q(net192));
 sky130_fd_sc_hd__dfxtp_4 _6913_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0048_),
    .Q(net193));
 sky130_fd_sc_hd__dfxtp_4 _6914_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0049_),
    .Q(net179));
 sky130_fd_sc_hd__dfxtp_4 _6915_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0050_),
    .Q(net180));
 sky130_fd_sc_hd__dfxtp_4 _6916_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0051_),
    .Q(net181));
 sky130_fd_sc_hd__dfxtp_4 _6917_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0052_),
    .Q(net182));
 sky130_fd_sc_hd__dfxtp_4 _6918_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0053_),
    .Q(net183));
 sky130_fd_sc_hd__dfxtp_4 _6919_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0054_),
    .Q(net184));
 sky130_fd_sc_hd__dfxtp_1 _6920_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0055_),
    .Q(\core_0.dec_mem_access ));
 sky130_fd_sc_hd__dfxtp_2 _6921_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0056_),
    .Q(\core_0.dec_mem_we ));
 sky130_fd_sc_hd__dfxtp_1 _6922_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0057_),
    .Q(\core_0.dec_used_operands[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6923_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0058_),
    .Q(\core_0.dec_used_operands[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6924_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0059_),
    .Q(\core_0.dec_sreg_load ));
 sky130_fd_sc_hd__dfxtp_2 _6925_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0060_),
    .Q(\core_0.dec_sreg_store ));
 sky130_fd_sc_hd__dfxtp_4 _6926_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0061_),
    .Q(\core_0.dec_sreg_jal_over ));
 sky130_fd_sc_hd__dfxtp_2 _6927_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0062_),
    .Q(\core_0.dec_sreg_irt ));
 sky130_fd_sc_hd__dfxtp_1 _6928_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0063_),
    .Q(\core_0.dec_sys ));
 sky130_fd_sc_hd__dfxtp_1 _6929_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0064_),
    .Q(\core_0.dec_mem_width ));
 sky130_fd_sc_hd__dfxtp_1 _6930_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0065_),
    .Q(\core_0.dec_mem_long ));
 sky130_fd_sc_hd__dfxtp_1 _6931_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0066_),
    .Q(\core_0.decode.input_valid ));
 sky130_fd_sc_hd__dfxtp_1 _6932_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0067_),
    .Q(\core_0.execute.sreg_priv_control.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6933_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0068_),
    .Q(\core_0.execute.sreg_data_page ));
 sky130_fd_sc_hd__dfxtp_2 _6934_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0069_),
    .Q(\core_0.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__dfxtp_1 _6935_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0070_),
    .Q(\core_0.execute.sreg_priv_control.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6936_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0071_),
    .Q(\core_0.execute.sreg_priv_control.o_d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6937_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0072_),
    .Q(\core_0.execute.sreg_priv_control.o_d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6938_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0073_),
    .Q(\core_0.execute.sreg_priv_control.o_d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6939_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0074_),
    .Q(\core_0.execute.sreg_priv_control.o_d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6940_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0075_),
    .Q(\core_0.execute.sreg_priv_control.o_d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6941_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0076_),
    .Q(\core_0.execute.sreg_priv_control.o_d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6942_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0077_),
    .Q(\core_0.execute.sreg_priv_control.o_d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6943_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0078_),
    .Q(\core_0.execute.sreg_priv_control.o_d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6944_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0079_),
    .Q(\core_0.execute.sreg_priv_control.o_d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6945_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0080_),
    .Q(\core_0.execute.sreg_priv_control.o_d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6946_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0081_),
    .Q(\core_0.execute.sreg_priv_control.o_d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6947_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0082_),
    .Q(\core_0.execute.alu_mul_div.comp ));
 sky130_fd_sc_hd__dfxtp_1 _6948_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0083_),
    .Q(\core_0.fetch.out_buffer_data_instr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6949_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0084_),
    .Q(\core_0.fetch.out_buffer_data_instr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6950_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0085_),
    .Q(\core_0.fetch.out_buffer_data_instr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6951_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0086_),
    .Q(\core_0.fetch.out_buffer_data_instr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6952_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0087_),
    .Q(\core_0.fetch.out_buffer_data_instr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6953_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0088_),
    .Q(\core_0.fetch.out_buffer_data_instr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6954_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0089_),
    .Q(\core_0.fetch.out_buffer_data_instr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6955_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0090_),
    .Q(\core_0.fetch.out_buffer_data_instr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6956_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0091_),
    .Q(\core_0.fetch.out_buffer_data_instr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6957_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0092_),
    .Q(\core_0.fetch.out_buffer_data_instr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6958_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0093_),
    .Q(\core_0.fetch.out_buffer_data_instr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6959_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0094_),
    .Q(\core_0.fetch.out_buffer_data_instr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6960_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0095_),
    .Q(\core_0.fetch.out_buffer_data_instr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6961_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0096_),
    .Q(\core_0.fetch.out_buffer_data_instr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6962_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0097_),
    .Q(\core_0.fetch.out_buffer_data_instr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6963_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0098_),
    .Q(\core_0.fetch.out_buffer_data_instr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6964_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0099_),
    .Q(\core_0.fetch.out_buffer_data_instr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _6965_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0100_),
    .Q(\core_0.fetch.out_buffer_data_instr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _6966_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0101_),
    .Q(\core_0.fetch.out_buffer_data_instr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _6967_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0102_),
    .Q(\core_0.fetch.out_buffer_data_instr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _6968_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0103_),
    .Q(\core_0.fetch.out_buffer_data_instr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _6969_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0104_),
    .Q(\core_0.fetch.out_buffer_data_instr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _6970_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0105_),
    .Q(\core_0.fetch.out_buffer_data_instr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _6971_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0106_),
    .Q(\core_0.fetch.out_buffer_data_instr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _6972_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0107_),
    .Q(\core_0.fetch.out_buffer_data_instr[24] ));
 sky130_fd_sc_hd__dfxtp_1 _6973_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0108_),
    .Q(\core_0.fetch.out_buffer_data_instr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _6974_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0109_),
    .Q(\core_0.fetch.out_buffer_data_instr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _6975_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0110_),
    .Q(\core_0.fetch.out_buffer_data_instr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _6976_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0111_),
    .Q(\core_0.fetch.out_buffer_data_instr[28] ));
 sky130_fd_sc_hd__dfxtp_1 _6977_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0112_),
    .Q(\core_0.fetch.out_buffer_data_instr[29] ));
 sky130_fd_sc_hd__dfxtp_1 _6978_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0113_),
    .Q(\core_0.fetch.out_buffer_data_instr[30] ));
 sky130_fd_sc_hd__dfxtp_1 _6979_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0114_),
    .Q(\core_0.fetch.out_buffer_data_instr[31] ));
 sky130_fd_sc_hd__dfxtp_2 _6980_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0115_),
    .Q(\core_0.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__dfxtp_1 _6981_ (.CLK(clknet_leaf_27_i_clk),
    .D(\core_0.fetch.current_req_branch_pred ),
    .Q(\core_0.fetch.prev_req_branch_pred ));
 sky130_fd_sc_hd__dfxtp_1 _6982_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0116_),
    .Q(\core_0.fetch.prev_request_pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6983_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0117_),
    .Q(\core_0.fetch.prev_request_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6984_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0118_),
    .Q(\core_0.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6985_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0119_),
    .Q(\core_0.fetch.prev_request_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6986_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0120_),
    .Q(\core_0.fetch.prev_request_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6987_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0121_),
    .Q(\core_0.fetch.prev_request_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6988_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0122_),
    .Q(\core_0.fetch.prev_request_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6989_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0123_),
    .Q(\core_0.fetch.prev_request_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6990_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0124_),
    .Q(\core_0.fetch.prev_request_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6991_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0125_),
    .Q(\core_0.fetch.prev_request_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6992_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0126_),
    .Q(\core_0.fetch.prev_request_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6993_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0127_),
    .Q(\core_0.fetch.prev_request_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6994_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0128_),
    .Q(\core_0.fetch.prev_request_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6995_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0129_),
    .Q(\core_0.fetch.prev_request_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6996_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0130_),
    .Q(\core_0.fetch.prev_request_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6997_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0131_),
    .Q(\core_0.fetch.prev_request_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6998_ (.CLK(clknet_leaf_28_i_clk),
    .D(\core_0.fetch.submitable ),
    .Q(\core_0.decode.i_submit ));
 sky130_fd_sc_hd__dfxtp_1 _6999_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0132_),
    .Q(\core_0.fetch.out_buffer_data_pred ));
 sky130_fd_sc_hd__dfxtp_4 _7000_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0133_),
    .Q(\core_0.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7001_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0134_),
    .Q(\core_0.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7002_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0135_),
    .Q(\core_0.decode.i_instr_l[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7003_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0136_),
    .Q(\core_0.decode.i_instr_l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7004_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0137_),
    .Q(\core_0.decode.i_instr_l[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7005_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0138_),
    .Q(\core_0.decode.i_instr_l[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7006_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0139_),
    .Q(\core_0.decode.i_instr_l[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7007_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0140_),
    .Q(\core_0.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7008_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0141_),
    .Q(\core_0.decode.i_instr_l[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7009_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0142_),
    .Q(\core_0.decode.i_instr_l[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7010_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0143_),
    .Q(\core_0.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7011_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0144_),
    .Q(\core_0.decode.i_instr_l[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7012_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0145_),
    .Q(\core_0.decode.i_instr_l[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7013_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0146_),
    .Q(\core_0.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7014_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0147_),
    .Q(\core_0.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7015_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0148_),
    .Q(\core_0.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7016_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0149_),
    .Q(\core_0.decode.i_imm_pass[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7017_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0150_),
    .Q(\core_0.decode.i_imm_pass[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7018_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0151_),
    .Q(\core_0.decode.i_imm_pass[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7019_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0152_),
    .Q(\core_0.decode.i_imm_pass[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7020_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0153_),
    .Q(\core_0.decode.i_imm_pass[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7021_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0154_),
    .Q(\core_0.decode.i_imm_pass[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7022_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0155_),
    .Q(\core_0.decode.i_imm_pass[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7023_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0156_),
    .Q(\core_0.decode.i_imm_pass[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7024_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0157_),
    .Q(\core_0.decode.i_imm_pass[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7025_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0158_),
    .Q(\core_0.decode.i_imm_pass[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7026_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0159_),
    .Q(\core_0.decode.i_imm_pass[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7027_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0160_),
    .Q(\core_0.decode.i_imm_pass[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7028_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0161_),
    .Q(\core_0.decode.i_imm_pass[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7029_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0162_),
    .Q(\core_0.decode.i_imm_pass[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7030_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0163_),
    .Q(\core_0.decode.i_imm_pass[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7031_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0164_),
    .Q(\core_0.decode.i_imm_pass[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7032_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0165_),
    .Q(\core_0.fetch.dbg_out ));
 sky130_fd_sc_hd__dfxtp_1 _7033_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0166_),
    .Q(\core_0.fetch.flush_event_invalidate ));
 sky130_fd_sc_hd__dfxtp_1 _7034_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0167_),
    .Q(\core_0.fetch.pc_flush_override ));
 sky130_fd_sc_hd__dfxtp_1 _7035_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0168_),
    .Q(\core_0.fetch.pc_reset_override ));
 sky130_fd_sc_hd__dfxtp_2 _7036_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0169_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _7037_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0170_),
    .Q(\core_0.decode.i_jmp_pred_pass ));
 sky130_fd_sc_hd__dfxtp_1 _7038_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0004_),
    .Q(\core_0.decode.oc_alu_mode[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7039_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0005_),
    .Q(\core_0.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7040_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0006_),
    .Q(\core_0.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__dfxtp_2 _7041_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0007_),
    .Q(\core_0.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7042_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0008_),
    .Q(\core_0.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__dfxtp_2 _7043_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0009_),
    .Q(\core_0.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7044_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0010_),
    .Q(\core_0.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__dfxtp_2 _7045_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0011_),
    .Q(\core_0.execute.alu_mul_div.i_mul ));
 sky130_fd_sc_hd__dfxtp_2 _7046_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0012_),
    .Q(\core_0.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__dfxtp_4 _7047_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0000_),
    .Q(\core_0.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__dfxtp_4 _7048_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0001_),
    .Q(\core_0.decode.oc_alu_mode[11] ));
 sky130_fd_sc_hd__dfxtp_4 _7049_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0002_),
    .Q(\core_0.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7050_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0003_),
    .Q(\core_0.decode.oc_alu_mode[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7051_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0171_),
    .Q(\core_0.execute.alu_mul_div.div_cur[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7052_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0172_),
    .Q(\core_0.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7053_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0173_),
    .Q(\core_0.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__dfxtp_2 _7054_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0174_),
    .Q(\core_0.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7055_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0175_),
    .Q(\core_0.execute.alu_mul_div.div_cur[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7056_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0176_),
    .Q(\core_0.execute.alu_mul_div.div_cur[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7057_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0177_),
    .Q(\core_0.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7058_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0178_),
    .Q(\core_0.execute.alu_mul_div.div_cur[8] ));
 sky130_fd_sc_hd__dfxtp_2 _7059_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0179_),
    .Q(\core_0.execute.alu_mul_div.div_cur[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7060_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0180_),
    .Q(\core_0.execute.alu_mul_div.div_cur[10] ));
 sky130_fd_sc_hd__dfxtp_2 _7061_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0181_),
    .Q(\core_0.execute.alu_mul_div.div_cur[11] ));
 sky130_fd_sc_hd__dfxtp_2 _7062_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0182_),
    .Q(\core_0.execute.alu_mul_div.div_cur[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7063_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0183_),
    .Q(\core_0.execute.alu_mul_div.div_cur[13] ));
 sky130_fd_sc_hd__dfxtp_2 _7064_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0184_),
    .Q(\core_0.execute.alu_mul_div.div_cur[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7065_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0185_),
    .Q(\core_0.execute.alu_mul_div.div_cur[15] ));
 sky130_fd_sc_hd__dfxtp_2 _7066_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0186_),
    .Q(\core_0.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__dfxtp_4 _7067_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0187_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_4 _7068_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0188_),
    .Q(\core_0.execute.alu_mul_div.cbit[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7069_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0189_),
    .Q(\core_0.execute.alu_mul_div.cbit[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7070_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0190_),
    .Q(\core_0.execute.alu_mul_div.cbit[3] ));
 sky130_fd_sc_hd__dfxtp_2 _7071_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0191_),
    .Q(\core_0.de_jmp_pred ));
 sky130_fd_sc_hd__dfxtp_1 _7072_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0192_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_1 _7073_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0014_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_1 _7074_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0193_),
    .Q(\core_0.execute.mem_stage_pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7075_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0194_),
    .Q(\core_0.execute.mem_stage_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7076_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0195_),
    .Q(\core_0.execute.mem_stage_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7077_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0196_),
    .Q(\core_0.execute.mem_stage_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7078_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0197_),
    .Q(\core_0.execute.mem_stage_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7079_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0198_),
    .Q(\core_0.execute.mem_stage_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7080_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0199_),
    .Q(\core_0.execute.mem_stage_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7081_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0200_),
    .Q(\core_0.execute.mem_stage_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7082_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0201_),
    .Q(\core_0.execute.mem_stage_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7083_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0202_),
    .Q(\core_0.execute.mem_stage_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7084_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0203_),
    .Q(\core_0.execute.mem_stage_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7085_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0204_),
    .Q(\core_0.execute.mem_stage_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7086_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0205_),
    .Q(\core_0.execute.mem_stage_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7087_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0206_),
    .Q(\core_0.execute.mem_stage_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7088_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0207_),
    .Q(\core_0.execute.mem_stage_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7089_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0208_),
    .Q(\core_0.execute.mem_stage_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7090_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0209_),
    .Q(\core_0.execute.prev_pc_high[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7091_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0210_),
    .Q(\core_0.execute.prev_pc_high[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7092_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0211_),
    .Q(\core_0.execute.prev_pc_high[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7093_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0212_),
    .Q(\core_0.execute.prev_pc_high[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7094_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0213_),
    .Q(\core_0.execute.prev_pc_high[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7095_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0214_),
    .Q(\core_0.execute.prev_pc_high[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7096_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0215_),
    .Q(\core_0.execute.prev_pc_high[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7097_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0216_),
    .Q(\core_0.execute.prev_pc_high[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7098_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0217_),
    .Q(\core_0.execute.sreg_irq_flags.i_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7099_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0218_),
    .Q(\core_0.execute.prev_sys ));
 sky130_fd_sc_hd__dfxtp_1 _7100_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0219_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_1 _7101_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0220_),
    .Q(\core_0.ew_addr_high[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7102_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0221_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_1 _7103_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0222_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_2 _7104_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0223_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_2 _7105_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0224_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_2 _7106_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0225_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_2 _7107_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0226_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_2 _7108_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0227_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_2 _7109_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0228_),
    .Q(\core_0.ew_submit ));
 sky130_fd_sc_hd__dfxtp_2 _7110_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0229_),
    .Q(\core_0.ew_data[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7111_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0230_),
    .Q(\core_0.ew_data[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7112_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0231_),
    .Q(\core_0.ew_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7113_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0232_),
    .Q(\core_0.ew_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7114_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0233_),
    .Q(\core_0.ew_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7115_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0234_),
    .Q(\core_0.ew_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7116_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0235_),
    .Q(\core_0.ew_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7117_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0236_),
    .Q(\core_0.ew_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7118_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0237_),
    .Q(\core_0.ew_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7119_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0238_),
    .Q(\core_0.ew_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7120_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0239_),
    .Q(\core_0.ew_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7121_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0240_),
    .Q(\core_0.ew_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7122_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0241_),
    .Q(\core_0.ew_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7123_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0242_),
    .Q(\core_0.ew_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7124_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0243_),
    .Q(\core_0.ew_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7125_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0244_),
    .Q(\core_0.ew_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7126_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0245_),
    .Q(\core_0.ew_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7127_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0246_),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_1 _7128_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0247_),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_1 _7129_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0248_),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_1 _7130_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0249_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_1 _7131_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0250_),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_1 _7132_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0251_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_1 _7133_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0252_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_1 _7134_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0253_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_1 _7135_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0254_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _7136_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0255_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_1 _7137_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0256_),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_1 _7138_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0257_),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_1 _7139_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0258_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_1 _7140_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0259_),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_1 _7141_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0260_),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_1 _7142_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0261_),
    .Q(\core_0.ew_reg_ie[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7143_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0262_),
    .Q(\core_0.ew_reg_ie[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7144_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0263_),
    .Q(\core_0.ew_reg_ie[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7145_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0264_),
    .Q(\core_0.ew_reg_ie[3] ));
 sky130_fd_sc_hd__dfxtp_4 _7146_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0265_),
    .Q(\core_0.ew_reg_ie[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7147_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0266_),
    .Q(\core_0.ew_reg_ie[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7148_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0267_),
    .Q(\core_0.ew_reg_ie[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7149_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0268_),
    .Q(\core_0.ew_reg_ie[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7150_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0269_),
    .Q(\core_0.ew_mem_access ));
 sky130_fd_sc_hd__dfxtp_2 _7151_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0270_),
    .Q(\core_0.ew_mem_width ));
 sky130_fd_sc_hd__dfxtp_1 _7152_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0013_),
    .Q(\core_0.decode.i_flush ));
 sky130_fd_sc_hd__dfxtp_2 _7153_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0271_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _7154_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0272_),
    .Q(\core_0.execute.hold_valid ));
 sky130_fd_sc_hd__dfxtp_1 _7155_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0273_),
    .Q(\core_0.execute.rf.reg_outputs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7156_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0274_),
    .Q(\core_0.execute.rf.reg_outputs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7157_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0275_),
    .Q(\core_0.execute.rf.reg_outputs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7158_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0276_),
    .Q(\core_0.execute.rf.reg_outputs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7159_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0277_),
    .Q(\core_0.execute.rf.reg_outputs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7160_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0278_),
    .Q(\core_0.execute.rf.reg_outputs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7161_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0279_),
    .Q(\core_0.execute.rf.reg_outputs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7162_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0280_),
    .Q(\core_0.execute.rf.reg_outputs[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7163_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0281_),
    .Q(\core_0.execute.rf.reg_outputs[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7164_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0282_),
    .Q(\core_0.execute.rf.reg_outputs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7165_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0283_),
    .Q(\core_0.execute.rf.reg_outputs[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7166_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0284_),
    .Q(\core_0.execute.rf.reg_outputs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7167_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0285_),
    .Q(\core_0.execute.rf.reg_outputs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7168_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0286_),
    .Q(\core_0.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7169_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0287_),
    .Q(\core_0.execute.rf.reg_outputs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7170_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0288_),
    .Q(\core_0.execute.rf.reg_outputs[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7171_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0289_),
    .Q(\core_0.execute.rf.reg_outputs[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7172_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0290_),
    .Q(\core_0.execute.rf.reg_outputs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7173_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0291_),
    .Q(\core_0.execute.rf.reg_outputs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7174_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0292_),
    .Q(\core_0.execute.rf.reg_outputs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7175_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0293_),
    .Q(\core_0.execute.rf.reg_outputs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7176_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0294_),
    .Q(\core_0.execute.rf.reg_outputs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7177_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0295_),
    .Q(\core_0.execute.rf.reg_outputs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7178_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0296_),
    .Q(\core_0.execute.rf.reg_outputs[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7179_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0297_),
    .Q(\core_0.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7180_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0298_),
    .Q(\core_0.execute.rf.reg_outputs[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7181_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0299_),
    .Q(\core_0.execute.rf.reg_outputs[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7182_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0300_),
    .Q(\core_0.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7183_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0301_),
    .Q(\core_0.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7184_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0302_),
    .Q(\core_0.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7185_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0303_),
    .Q(\core_0.execute.rf.reg_outputs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7186_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0304_),
    .Q(\core_0.execute.rf.reg_outputs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7187_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0305_),
    .Q(\core_0.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7188_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0306_),
    .Q(\core_0.execute.rf.reg_outputs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7189_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0307_),
    .Q(\core_0.execute.rf.reg_outputs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7190_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0308_),
    .Q(\core_0.execute.rf.reg_outputs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7191_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0309_),
    .Q(\core_0.execute.rf.reg_outputs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7192_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0310_),
    .Q(\core_0.execute.rf.reg_outputs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7193_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0311_),
    .Q(\core_0.execute.rf.reg_outputs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7194_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0312_),
    .Q(\core_0.execute.rf.reg_outputs[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7195_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0313_),
    .Q(\core_0.execute.rf.reg_outputs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7196_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0314_),
    .Q(\core_0.execute.rf.reg_outputs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7197_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0315_),
    .Q(\core_0.execute.rf.reg_outputs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7198_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0316_),
    .Q(\core_0.execute.rf.reg_outputs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7199_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0317_),
    .Q(\core_0.execute.rf.reg_outputs[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7200_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0318_),
    .Q(\core_0.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7201_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0319_),
    .Q(\core_0.execute.rf.reg_outputs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7202_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0320_),
    .Q(\core_0.execute.rf.reg_outputs[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _7203_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0321_),
    .Q(\core_0.execute.rf.reg_outputs[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _7204_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0322_),
    .Q(\core_0.execute.rf.reg_outputs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7205_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0323_),
    .Q(\core_0.execute.rf.reg_outputs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7206_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0324_),
    .Q(\core_0.execute.rf.reg_outputs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7207_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0325_),
    .Q(\core_0.execute.rf.reg_outputs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7208_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0326_),
    .Q(\core_0.execute.rf.reg_outputs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7209_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0327_),
    .Q(\core_0.execute.rf.reg_outputs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7210_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0328_),
    .Q(\core_0.execute.rf.reg_outputs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7211_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0329_),
    .Q(\core_0.execute.rf.reg_outputs[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7212_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0330_),
    .Q(\core_0.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7213_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0331_),
    .Q(\core_0.execute.rf.reg_outputs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7214_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0332_),
    .Q(\core_0.execute.rf.reg_outputs[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _7215_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0333_),
    .Q(\core_0.execute.rf.reg_outputs[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7216_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0334_),
    .Q(\core_0.execute.rf.reg_outputs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7217_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0335_),
    .Q(\core_0.execute.rf.reg_outputs[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7218_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0336_),
    .Q(\core_0.execute.rf.reg_outputs[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _7219_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0337_),
    .Q(\core_0.execute.rf.reg_outputs[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _7220_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0338_),
    .Q(\core_0.execute.rf.reg_outputs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7221_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0339_),
    .Q(\core_0.execute.rf.reg_outputs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7222_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0340_),
    .Q(\core_0.execute.rf.reg_outputs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7223_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0341_),
    .Q(\core_0.execute.rf.reg_outputs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7224_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0342_),
    .Q(\core_0.execute.rf.reg_outputs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7225_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0343_),
    .Q(\core_0.execute.rf.reg_outputs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7226_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0344_),
    .Q(\core_0.execute.rf.reg_outputs[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7227_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0345_),
    .Q(\core_0.execute.rf.reg_outputs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7228_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0346_),
    .Q(\core_0.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7229_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0347_),
    .Q(\core_0.execute.rf.reg_outputs[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7230_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0348_),
    .Q(\core_0.execute.rf.reg_outputs[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7231_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0349_),
    .Q(\core_0.execute.rf.reg_outputs[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _7232_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0350_),
    .Q(\core_0.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7233_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0351_),
    .Q(\core_0.execute.rf.reg_outputs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7234_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0352_),
    .Q(\core_0.execute.rf.reg_outputs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7235_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0353_),
    .Q(\core_0.execute.rf.reg_outputs[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7236_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0354_),
    .Q(\core_0.execute.rf.reg_outputs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7237_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0355_),
    .Q(\core_0.execute.rf.reg_outputs[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7238_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0356_),
    .Q(\core_0.execute.rf.reg_outputs[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7239_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0357_),
    .Q(\core_0.execute.rf.reg_outputs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7240_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0358_),
    .Q(\core_0.execute.rf.reg_outputs[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7241_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0359_),
    .Q(\core_0.execute.rf.reg_outputs[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7242_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0360_),
    .Q(\core_0.execute.rf.reg_outputs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7243_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0361_),
    .Q(\core_0.execute.rf.reg_outputs[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7244_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0362_),
    .Q(\core_0.execute.rf.reg_outputs[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7245_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0363_),
    .Q(\core_0.execute.rf.reg_outputs[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7246_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0364_),
    .Q(\core_0.execute.rf.reg_outputs[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7247_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0365_),
    .Q(\core_0.execute.rf.reg_outputs[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7248_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0366_),
    .Q(\core_0.execute.rf.reg_outputs[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7249_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0367_),
    .Q(\core_0.execute.rf.reg_outputs[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7250_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0368_),
    .Q(\core_0.execute.rf.reg_outputs[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7251_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0369_),
    .Q(\core_0.execute.rf.reg_outputs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7252_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0370_),
    .Q(\core_0.execute.rf.reg_outputs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7253_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0371_),
    .Q(\core_0.execute.rf.reg_outputs[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7254_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0372_),
    .Q(\core_0.execute.rf.reg_outputs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7255_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0373_),
    .Q(\core_0.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7256_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0374_),
    .Q(\core_0.execute.rf.reg_outputs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7257_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0375_),
    .Q(\core_0.execute.rf.reg_outputs[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _7258_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0376_),
    .Q(\core_0.execute.rf.reg_outputs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7259_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0377_),
    .Q(\core_0.execute.rf.reg_outputs[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7260_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0378_),
    .Q(\core_0.execute.rf.reg_outputs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7261_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0379_),
    .Q(\core_0.execute.rf.reg_outputs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7262_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0380_),
    .Q(\core_0.execute.rf.reg_outputs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7263_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0381_),
    .Q(\core_0.execute.rf.reg_outputs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7264_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0382_),
    .Q(\core_0.execute.rf.reg_outputs[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7265_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0383_),
    .Q(\core_0.execute.rf.reg_outputs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7266_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0384_),
    .Q(\core_0.execute.rf.reg_outputs[1][15] ));
 sky130_fd_sc_hd__dfxtp_4 _7267_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0385_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_4 _7268_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0386_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_4 _7269_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0387_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_4 _7270_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0388_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_4 _7271_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0389_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_4 _7272_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0390_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_4 _7273_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0391_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_4 _7274_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0392_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_4 _7275_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0393_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_4 _7276_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0394_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_4 _7277_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0395_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_4 _7278_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0396_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_4 _7279_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0397_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_4 _7280_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0398_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_4 _7281_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0399_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_2 _7282_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0400_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_1 _7283_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0401_),
    .Q(\core_0.execute.irq_en ));
 sky130_fd_sc_hd__dfxtp_2 _7284_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0402_),
    .Q(\core_0.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7285_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0403_),
    .Q(\core_0.execute.alu_mul_div.mul_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7286_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0404_),
    .Q(\core_0.execute.alu_mul_div.mul_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7287_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0405_),
    .Q(\core_0.execute.alu_mul_div.mul_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7288_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0406_),
    .Q(\core_0.execute.alu_mul_div.mul_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7289_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0407_),
    .Q(\core_0.execute.alu_mul_div.mul_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7290_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0408_),
    .Q(\core_0.execute.alu_mul_div.mul_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7291_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0409_),
    .Q(\core_0.execute.alu_mul_div.mul_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7292_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0410_),
    .Q(\core_0.execute.alu_mul_div.mul_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7293_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0411_),
    .Q(\core_0.execute.alu_mul_div.mul_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7294_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0412_),
    .Q(\core_0.execute.alu_mul_div.mul_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7295_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0413_),
    .Q(\core_0.execute.alu_mul_div.mul_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7296_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0414_),
    .Q(\core_0.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__dfxtp_2 _7297_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0415_),
    .Q(\core_0.execute.alu_mul_div.mul_res[12] ));
 sky130_fd_sc_hd__dfxtp_2 _7298_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0416_),
    .Q(\core_0.execute.alu_mul_div.mul_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7299_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0417_),
    .Q(\core_0.execute.alu_mul_div.mul_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7300_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0418_),
    .Q(\core_0.execute.alu_mul_div.mul_res[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7301_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0419_),
    .Q(\core_0.execute.next_ready_delayed ));
 sky130_fd_sc_hd__dfxtp_1 _7302_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0420_),
    .Q(\core_0.execute.alu_mul_div.div_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7303_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0421_),
    .Q(\core_0.execute.alu_mul_div.div_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7304_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0422_),
    .Q(\core_0.execute.alu_mul_div.div_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7305_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0423_),
    .Q(\core_0.execute.alu_mul_div.div_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7306_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0424_),
    .Q(\core_0.execute.alu_mul_div.div_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7307_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0425_),
    .Q(\core_0.execute.alu_mul_div.div_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7308_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0426_),
    .Q(\core_0.execute.alu_mul_div.div_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7309_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0427_),
    .Q(\core_0.execute.alu_mul_div.div_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7310_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0428_),
    .Q(\core_0.execute.alu_mul_div.div_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7311_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0429_),
    .Q(\core_0.execute.alu_mul_div.div_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7312_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0430_),
    .Q(\core_0.execute.alu_mul_div.div_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7313_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0431_),
    .Q(\core_0.execute.alu_mul_div.div_res[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7314_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0432_),
    .Q(\core_0.execute.alu_mul_div.div_res[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7315_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0433_),
    .Q(\core_0.execute.alu_mul_div.div_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7316_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0434_),
    .Q(\core_0.execute.alu_mul_div.div_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7317_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0435_),
    .Q(\core_0.execute.alu_mul_div.div_res[15] ));
 sky130_fd_sc_hd__dfxtp_4 _7318_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0436_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_4 _7319_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0437_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_4 _7320_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0438_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_4 _7321_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0439_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_4 _7322_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0440_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_4 _7323_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0441_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_4 _7324_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0442_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_4 _7325_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0443_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_4 _7326_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0444_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_4 _7327_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0445_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_4 _7328_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0446_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_4 _7329_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0447_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_4 _7330_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0448_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_4 _7331_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0449_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_4 _7332_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0450_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_2 _7333_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0451_),
    .Q(\core_0.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_4 _7334_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0452_),
    .Q(\core_0.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7335_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0453_),
    .Q(\core_0.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7336_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0454_),
    .Q(\core_0.execute.alu_flag_reg.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7337_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0455_),
    .Q(\core_0.execute.alu_flag_reg.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7338_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0456_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7339_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0457_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7340_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0458_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7341_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0459_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7342_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0460_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7343_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0461_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7344_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0462_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7345_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0463_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[7] ));
 sky130_fd_sc_hd__dfxtp_2 _7346_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0464_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7347_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0465_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7348_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0466_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7349_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0467_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7350_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0468_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7351_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0469_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7352_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0470_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7353_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0471_),
    .Q(\core_0.execute.sreg_irq_pc.o_d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7354_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0472_),
    .Q(\core_0.execute.sreg_jtr_buff.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7355_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0473_),
    .Q(\core_0.execute.sreg_jtr_buff.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7356_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0474_),
    .Q(\core_0.execute.sreg_jtr_buff.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7357_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0475_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_1 _7358_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0476_),
    .Q(\core_0.execute.trap_flag ));
 sky130_fd_sc_hd__dfxtp_4 _7359_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0477_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_1 _7360_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0478_),
    .Q(\core_0.execute.sreg_scratch.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7361_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0479_),
    .Q(\core_0.execute.sreg_scratch.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7362_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0480_),
    .Q(\core_0.execute.sreg_scratch.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7363_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0481_),
    .Q(\core_0.execute.sreg_scratch.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7364_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0482_),
    .Q(\core_0.execute.sreg_scratch.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7365_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0483_),
    .Q(\core_0.execute.sreg_scratch.o_d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7366_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0484_),
    .Q(\core_0.execute.sreg_scratch.o_d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7367_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0485_),
    .Q(\core_0.execute.sreg_scratch.o_d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7368_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0486_),
    .Q(\core_0.execute.sreg_scratch.o_d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7369_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0487_),
    .Q(\core_0.execute.sreg_scratch.o_d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7370_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0488_),
    .Q(\core_0.execute.sreg_scratch.o_d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7371_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0489_),
    .Q(\core_0.execute.sreg_scratch.o_d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7372_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0490_),
    .Q(\core_0.execute.sreg_scratch.o_d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7373_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0491_),
    .Q(\core_0.execute.sreg_scratch.o_d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7374_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0492_),
    .Q(\core_0.execute.sreg_scratch.o_d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7375_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0493_),
    .Q(\core_0.execute.sreg_scratch.o_d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7376_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0494_),
    .Q(\core_0.execute.sreg_irq_flags.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7377_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0495_),
    .Q(\core_0.execute.sreg_irq_flags.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7378_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0496_),
    .Q(\core_0.execute.sreg_irq_flags.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7379_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0497_),
    .Q(\core_0.execute.sreg_irq_flags.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7380_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0498_),
    .Q(\core_0.execute.sreg_irq_flags.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7381_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0499_),
    .Q(\core_0.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7382_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0500_),
    .Q(\core_0.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7383_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0501_),
    .Q(\core_0.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7384_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0502_),
    .Q(\core_0.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__dfxtp_2 _7385_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0503_),
    .Q(\core_0.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7386_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0504_),
    .Q(\core_0.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7387_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0505_),
    .Q(\core_0.execute.pc_high_out[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7388_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0506_),
    .Q(\core_0.execute.pc_high_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7389_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0507_),
    .Q(\core_0.execute.pc_high_buff_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7390_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0508_),
    .Q(\core_0.execute.pc_high_buff_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7391_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0509_),
    .Q(\core_0.execute.pc_high_buff_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7392_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0510_),
    .Q(\core_0.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7393_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0511_),
    .Q(\core_0.execute.pc_high_buff_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7394_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0512_),
    .Q(\core_0.execute.pc_high_buff_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7395_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0513_),
    .Q(\core_0.execute.pc_high_buff_out[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7396_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0514_),
    .Q(\core_0.execute.pc_high_buff_out[7] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(i_core_int_sreg[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(i_core_int_sreg[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(i_core_int_sreg[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(i_core_int_sreg[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(i_core_int_sreg[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(i_core_int_sreg[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(i_core_int_sreg[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(i_core_int_sreg[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(i_core_int_sreg[2]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(i_core_int_sreg[3]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(i_core_int_sreg[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(i_core_int_sreg[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(i_core_int_sreg[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(i_core_int_sreg[7]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(i_core_int_sreg[8]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(i_core_int_sreg[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(i_disable),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(i_irq),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(i_mc_core_int),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(i_mem_ack),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(i_mem_data[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(i_mem_data[10]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(i_mem_data[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(i_mem_data[12]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(i_mem_data[13]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(i_mem_data[14]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(i_mem_data[15]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(i_mem_data[1]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(i_mem_data[2]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(i_mem_data[3]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(i_mem_data[4]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(i_mem_data[5]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(i_mem_data[6]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(i_mem_data[7]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(i_mem_data[8]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(i_mem_data[9]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(i_mem_exception),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(i_req_data[0]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(i_req_data[10]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(i_req_data[11]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(i_req_data[12]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(i_req_data[13]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(i_req_data[14]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(i_req_data[15]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(i_req_data[16]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(i_req_data[17]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(i_req_data[18]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(i_req_data[19]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 input49 (.A(i_req_data[1]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(i_req_data[20]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(i_req_data[21]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(i_req_data[22]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(i_req_data[23]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(i_req_data[24]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(i_req_data[25]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(i_req_data[26]),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(i_req_data[27]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(i_req_data[28]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(i_req_data[29]),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input60 (.A(i_req_data[2]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(i_req_data[30]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(i_req_data[31]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(i_req_data[3]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(i_req_data[4]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(i_req_data[5]),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(i_req_data[6]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(i_req_data[7]),
    .X(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 input68 (.A(i_req_data[8]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(i_req_data[9]),
    .X(net69));
 sky130_fd_sc_hd__buf_6 input70 (.A(i_req_data_valid),
    .X(net70));
 sky130_fd_sc_hd__buf_6 input71 (.A(i_rst),
    .X(net71));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(dbg_pc[0]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(dbg_pc[10]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(dbg_pc[11]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(dbg_pc[12]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(dbg_pc[13]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(dbg_pc[14]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(dbg_pc[15]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(dbg_pc[1]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(dbg_pc[2]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(dbg_pc[3]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(dbg_pc[4]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(dbg_pc[5]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(dbg_pc[6]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(dbg_pc[7]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(dbg_pc[8]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(dbg_pc[9]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(dbg_r0[0]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(dbg_r0[10]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(dbg_r0[11]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(dbg_r0[12]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(dbg_r0[13]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(dbg_r0[14]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(dbg_r0[15]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(dbg_r0[1]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(dbg_r0[2]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(dbg_r0[3]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(dbg_r0[4]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(dbg_r0[5]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(dbg_r0[6]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(dbg_r0[7]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(dbg_r0[8]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(dbg_r0[9]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(o_c_data_page));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(o_c_instr_long));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(o_c_instr_page));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(o_icache_flush));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(o_instr_long_addr[0]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(o_instr_long_addr[1]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(o_instr_long_addr[2]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(o_instr_long_addr[3]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(o_instr_long_addr[4]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(o_instr_long_addr[5]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(o_instr_long_addr[6]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(o_instr_long_addr[7]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(o_mem_addr[0]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(o_mem_addr[10]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(o_mem_addr[11]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(o_mem_addr[12]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(o_mem_addr[13]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(o_mem_addr[14]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(o_mem_addr[15]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(o_mem_addr[1]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(o_mem_addr[2]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(o_mem_addr[3]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(o_mem_addr[4]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(o_mem_addr[5]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(o_mem_addr[6]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(o_mem_addr[7]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(o_mem_addr[8]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(o_mem_addr[9]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(o_mem_addr_high[0]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(o_mem_addr_high[1]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(o_mem_addr_high[2]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(o_mem_addr_high[3]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(o_mem_addr_high[4]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(o_mem_addr_high[5]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(o_mem_addr_high[6]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(o_mem_data[0]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(o_mem_data[10]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(o_mem_data[11]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(o_mem_data[12]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(o_mem_data[13]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(o_mem_data[14]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(o_mem_data[15]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(o_mem_data[1]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(o_mem_data[2]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(o_mem_data[3]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(o_mem_data[4]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(o_mem_data[5]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(o_mem_data[6]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(o_mem_data[7]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(o_mem_data[8]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(o_mem_data[9]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(o_mem_long));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(o_mem_req));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(o_mem_sel[0]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(o_mem_sel[1]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(o_mem_we));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(o_req_active));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(o_req_addr[0]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(o_req_addr[10]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(o_req_addr[11]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(o_req_addr[12]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(o_req_addr[13]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(o_req_addr[14]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(o_req_addr[15]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(o_req_addr[1]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(o_req_addr[2]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(o_req_addr[3]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(o_req_addr[4]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(o_req_addr[5]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(o_req_addr[6]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(o_req_addr[7]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(o_req_addr[8]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(o_req_addr[9]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(o_req_ppl_submit));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(sr_bus_addr[0]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(sr_bus_addr[10]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(sr_bus_addr[11]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(sr_bus_addr[12]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(sr_bus_addr[13]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(sr_bus_addr[14]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(sr_bus_addr[15]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(sr_bus_addr[1]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(sr_bus_addr[2]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(sr_bus_addr[3]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(sr_bus_addr[4]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(sr_bus_addr[5]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(sr_bus_addr[6]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(sr_bus_addr[7]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(sr_bus_addr[8]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(sr_bus_addr[9]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(sr_bus_data_o[0]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(sr_bus_data_o[10]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(sr_bus_data_o[11]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(sr_bus_data_o[12]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(sr_bus_data_o[13]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(sr_bus_data_o[14]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(sr_bus_data_o[15]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(sr_bus_data_o[1]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(sr_bus_data_o[2]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(sr_bus_data_o[3]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(sr_bus_data_o[4]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(sr_bus_data_o[5]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(sr_bus_data_o[6]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(sr_bus_data_o[7]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(sr_bus_data_o[8]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(sr_bus_data_o[9]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(sr_bus_we));
 sky130_fd_sc_hd__conb_1 core0_211 (.LO(net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_48_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_i_clk (.A(clknet_opt_1_1_i_clk),
    .X(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_i_clk (.A(clknet_1_0_0_i_clk),
    .X(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_i_clk (.A(clknet_1_1_0_i_clk),
    .X(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_opt_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_1_i_clk (.A(clknet_opt_1_0_i_clk),
    .X(clknet_opt_1_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__D (.DIODE(_0011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__D (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__D (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7301__D (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__B (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__B (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__A (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__B (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__B1 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__B1 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__B1 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__B1 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__B2 (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__B2 (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A2 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__B1 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A2 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A2 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__B1 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A2 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A2 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A2 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A2 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__B1 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A_N (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__B (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A_N (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__B (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A_N (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__B (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__C (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__D (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__C (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__B_N (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__B1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A2 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A2 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__B1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__B1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__B1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A2 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__B1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__B1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A2 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A2 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__C (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__A_N (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__B (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__C (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__A_N (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A_N (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__B (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A_N (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__D (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__A_N (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__B (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__B_N (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A_N (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__B (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__B (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__A_N (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__B_N (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__C (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__B (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__B_N (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__A_N (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__C (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__C (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__C (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A_N (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__C (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__D (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__C (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__B (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__C (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__B1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__S1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__S1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A_N (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__C (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__B (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__C (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__B (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__B_N (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A_N (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__S0 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__S0 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__B (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__D (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__C (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__B_N (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__A_N (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__C (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A_N (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A1 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A1 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__A (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__D (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__B (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A_N (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__A_N (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__C (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A_N (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A_N (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__B2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__B2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A2 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__B (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__B1 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__B1 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__B1 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__B1 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__B1 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__B1 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__A1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A2 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A2 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__A1 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__A (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__A0 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__A0 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__A0 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__A0 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__A (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A2 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A2 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A0 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__A (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__A1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__A (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A2 (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__A0 (.DIODE(_0655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__A1 (.DIODE(_0655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__A1 (.DIODE(_0655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A (.DIODE(_0655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A0 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__S (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__S (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__S (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A1 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__S (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__S (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__S (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__S (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__S (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__S (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__S (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__S (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__S (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__S (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__S (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__S (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__B1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__B (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__B1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__B (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__C1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__B (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__A2 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__B (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__A (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__B1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A2_N (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__B (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__A2_N (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__B1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__A1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__B (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A2 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A2_N (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__B (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__B1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__B1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__B (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__B (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__A1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__B1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A2_N (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A1 (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__C1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__B (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__D (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__D (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__D (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__D (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__D (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__D (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__D (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__D (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__D (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__B (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__A2 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__A2 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__C (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__D (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A_N (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__B (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__C (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A_N (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__C (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__C (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__C (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__A_N (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__B1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__A_N (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__B_N (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__B_N (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A_N (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__C (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__C (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A2 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A2 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__A2 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__A2 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__A1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__B (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A2 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__A2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__A (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__B_N (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__B_N (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__A_N (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A_N (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__C1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__B1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__C (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__C (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__B (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A_N (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__C (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__B (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__B (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__B (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__B (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__B2 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__B2 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__B2 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A3 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__A2 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__B2 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__B (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A2 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__C (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__B (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__B (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__A2 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A2 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__A (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__A2 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A2 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A2 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__A2 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__A (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A2 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A2 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__A2 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B2 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B2 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__B2 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A2 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__S (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__S (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__S0 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__B (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__B2 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A2 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__B (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__A2 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__A2 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A2 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__A2 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__C1 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A0 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__B1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A_N (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__B2 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__B (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__S (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__B (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__B (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__B1_N (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__B1_N (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__B1_N (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__B1_N (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__B1_N (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__B1_N (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__A (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__B (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A2 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__C1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__A1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__B1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__B1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__A1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__B1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__A (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__B (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__B (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__C (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__A (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__C (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__B (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__B (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__B (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__B (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__B (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__C (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__B (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__B1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__B1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A0 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A0 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__D_N (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A0 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__D_N (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__B_N (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__A0 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__A2 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__B1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A0 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__B (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__A0 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A2 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__B1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__C (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__A0 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__B1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A2 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__D (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A0 (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A1 (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A2 (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A2 (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__A0 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A1 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A2 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A1_N (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__B (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A0 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__B1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__B1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__C (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__A0 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__D (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A0 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A1 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A2 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__A2 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__A0 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__C (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A0 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A1 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__B1 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__B1 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__D (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A0 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A1 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A2 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A2 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__A (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A0 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__B (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__A0 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__B1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__B1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__D (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__C (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__A0 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__D_N (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__B (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__C (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__C (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__C (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__B (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__C (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__B (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__B (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__A (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__A (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__B (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__B (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A2 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A2 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A2 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A2 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A2 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A2 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A2 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A2 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A2 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A2 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A2_N (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__B (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A2_N (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A0 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A2 (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__S (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A2 (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A2 (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__S (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__A2 (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__S (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A2 (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__B1 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__B1 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B1 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__B1 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__B1 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__B1 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__B1 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__B (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__C1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__C1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__C1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__C1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__C1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__C1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__C1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__C1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__C1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__C1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__B (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__A (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__B (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__B (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__B (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__A (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__B (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__A (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__B (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__C (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__B (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__B (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__B (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A2 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A2 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__B1 (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__B1 (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__B1 (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__B1 (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__B1 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__B1 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A2 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A2 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A2 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A2 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A2 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A2 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A2 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A2 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__S (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__S (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__S (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__S (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__S (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__S (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__S (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A_N (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A1 (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A_N (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__A (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__B1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__C (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A2 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__B1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__A (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A_N (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__A_N (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__D (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__B2 (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__B (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A1 (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__B (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__B (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__B (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A2 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A1 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A2 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__B (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A3 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__B (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__B1 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__B1 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__B1 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A1 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__B1 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__B1 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__B1 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__B1 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A2 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A2 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__A2 (.DIODE(_0954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__A2 (.DIODE(_0954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__A2 (.DIODE(_0954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__A2 (.DIODE(_0954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A2 (.DIODE(_0954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__A2 (.DIODE(_0954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A2 (.DIODE(_0954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__B1 (.DIODE(_0954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__B1 (.DIODE(_0954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__B1 (.DIODE(_0954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__C1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__B (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__B1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__B2 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A2 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A2_N (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A2 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A2 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A2 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__A2 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A2 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A2 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A2 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A1 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__C (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__B2 (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__B1 (.DIODE(_0962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__C (.DIODE(_0962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A (.DIODE(_0962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__C (.DIODE(_0962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A1 (.DIODE(_0962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__B1 (.DIODE(_0962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A1 (.DIODE(_0962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__B2 (.DIODE(_0962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__C1 (.DIODE(_0962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A1 (.DIODE(_0962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A1 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A1 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A1 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__B2 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A1 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A1 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A1 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A1 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A1 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A1 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B2 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__B1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__B1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__B1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__C1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__B1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__B1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__B1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__B1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__B1_N (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A_N (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A2 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__B1 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__C1 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__B1 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__C1 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__C1 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__C1 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__A2 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__B2 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__B (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__C (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__B (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__A (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__B1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__C1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__C1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__C1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__C1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__C1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__C1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__B1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__C1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A1 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A1 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__B2 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A1 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__B2 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__B2 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__B2 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A1 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A1 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A1 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__S (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__S (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__S (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__S (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__S (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__S (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A (.DIODE(_1023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__S (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__S (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__A (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__B1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__C_N (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A2 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__B (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__B (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__B (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__B (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__B (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__A2 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A2 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A2 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A2 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__A2 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A2 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A2 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__A2 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A2 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__A1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__B (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__B (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__B (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__C (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__C (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__C (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__C (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__D (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__C (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__B (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__B (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__D (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__B (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A2 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A2 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__B (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A2 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A2 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A2 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A2 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__B (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__B (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__B (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__B1 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__B (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__B (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A2 (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__A2 (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A2 (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__B (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__C (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A2 (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__B (.DIODE(_1045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A (.DIODE(_1045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__B (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__B (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__B (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__B (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__B (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__B (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__B (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__B (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__B (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__B (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__C (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__C (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__C (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__C (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__C (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__C (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__C (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__C (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__C (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__C (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__B (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__B1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__B (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__C (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__C (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__B (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__C (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A2_N (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B1 (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__A3 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__A2 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A2 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A3 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__B1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__B1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__B1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__B2 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__C1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__D1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A1 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__B1 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__B1 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A1 (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__B (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__A2 (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A2 (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A2 (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__B1 (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__B1 (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__B1 (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A1 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__A2 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A2 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A2 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A2 (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A2 (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__B1 (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__B1 (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__B1 (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__A2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__A2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__D (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__C (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__B (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__B1 (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__B (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A1_N (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A1_N (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A0 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A1 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A1 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__B1 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A1 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__C1 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A1 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__B1 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A1 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__B1_N (.DIODE(_1149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A3 (.DIODE(_1149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__A (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__B1 (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__A (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__A (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__B (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__B (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__B (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__B (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__B (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__A1 (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A2 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A2 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A2 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__A2 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A2 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A2 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A2 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A1 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__B2 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A (.DIODE(_1157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__B1 (.DIODE(_1157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__C1 (.DIODE(_1157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__C1 (.DIODE(_1157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A (.DIODE(_1157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A (.DIODE(_1157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A (.DIODE(_1157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A (.DIODE(_1157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__B (.DIODE(_1157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__B (.DIODE(_1157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__B (.DIODE(_1158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__C (.DIODE(_1158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__B (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__A2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__A2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__A2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__A2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__B (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__A (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__A2 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__B1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__B1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__A (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__B1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__B1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__B1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__B1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__B1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__B1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__A (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__A (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A1 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__C1 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A1 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__A1 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A1 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__A (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__S1 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A2 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__A1 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__S (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__C1 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__A (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__S (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__S (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__S1 (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__S0 (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__S1 (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A1 (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__A1 (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__S (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__S (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__A (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__S1 (.DIODE(_1206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__S0 (.DIODE(_1206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__S (.DIODE(_1206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__S1 (.DIODE(_1206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A2 (.DIODE(_1206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__S (.DIODE(_1206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__S (.DIODE(_1206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A1_N (.DIODE(_1206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__S (.DIODE(_1206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A (.DIODE(_1206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A1 (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__S1 (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__S0 (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6237__B (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__A1 (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__A1 (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__B (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__B (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__B (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__B (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__A (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A1 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__A1 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__A (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A1 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A1 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A2 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__A2 (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A2 (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__D_N (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__B1 (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__S (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__S (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__S (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__A (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__S (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__S (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__S (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__S (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__S (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__S (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__S (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__S (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__S (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__S (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__S (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__S (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__S (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__S (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__S (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__S (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__S (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__S (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__S (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__S (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__S (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__S (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__S (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__S (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__S (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__S (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__S (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__S (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__S (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__S (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A_N (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__C (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__C (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__C (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__C (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__C (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__C (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__C (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__C (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__C (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__S (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__S (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__S (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__S (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__S (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__S (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__S (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__S (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__S (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__S (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__A1 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__S (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__S (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__S (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__S (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__S (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__S (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__S (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__S (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__B2 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__B2 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__B2 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__B2 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__B2 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__B2 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__B2 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__B2 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A1 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A1 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__B (.DIODE(_1325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__B (.DIODE(_1325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__B (.DIODE(_1325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__B (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__B (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__S (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__C1 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__A (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__C1 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__C1 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__S (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__C1 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__C1 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__C1 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__D (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__B (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__B2 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__A2 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__B (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__B (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__A (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A2 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__B1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__B1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__B1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__B (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__B (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__D1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A1 (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A2 (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A1 (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__A1 (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A1 (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A1 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A1 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__S (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__S (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__S (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__S (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A1 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__A (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__S (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__S (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A2 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__A1 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A2 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__B (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__A (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A2 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__A (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__B1 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__B (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__B (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__B1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__B1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__B1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__B (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__B (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__D1 (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__B (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__B2 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A2 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__B (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A_N (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__A (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A1 (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A1 (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__B1 (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__B (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__B (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__B (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__B (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__B (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__A (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__C1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__C1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__C1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__A1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__B (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__B (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__B (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A1 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__C (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A1 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A2 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__B (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__D (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A2 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__A (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__A (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__B (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__A1 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__B (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__B (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__B (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__C (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__A2 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A2 (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__D (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__B (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__D (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A2 (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A1 (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__B (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__B (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__A (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__B1 (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__A2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__B (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__S (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__S (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__S (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__S (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__S (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__S (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A2 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__A (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__C1 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__S (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__S (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__S (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__S (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__S (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__S (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__S (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__S (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__B1_N (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__B1_N (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__B1_N (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__B1_N (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__B1_N (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__B1_N (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__B1_N (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__B1_N (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A2 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__B (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A2 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A2 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A2 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A2 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A2 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A2 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__B1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__S0 (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__B1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__S0 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__S1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__S (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__S (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A1 (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__S (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__S (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__S (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__S (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__S1 (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A1 (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__S (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__B (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__B (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__B1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__B1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__B1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__B1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__C1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__C1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__C1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__C1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__C1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__C1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A1 (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__A (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A1 (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A1 (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__D1 (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__B1 (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__S (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__B (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__B1 (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__A1 (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__A (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A1 (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A1 (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A2 (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__C1 (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A1 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__A1 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__A1 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A1 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__A1 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A1 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__C1 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__C1 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__B (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__A (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__C1 (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__C1 (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__C1 (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__C1 (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__C1 (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__C1 (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__C1 (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__C1 (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__C1 (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A2 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__C (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A1 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__C (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__B (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A2 (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A1 (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__A (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__B (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__B (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A0 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__A1 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A1 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__B1 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__B1 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__B1 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A2 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__B1 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__B1 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__A2 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A2 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A2 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A2 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__B1 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__C (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A2 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__A (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A2 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A2 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A2 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A2 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__A3 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A3 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A3 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A3 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A3 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__A3 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__B1 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__B1 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A2 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__A2 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__A2 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__A2 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A2 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__A2 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__B (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__B (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__A_N (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__A (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__A (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__D_N (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__A (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__C (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__A (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__C (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__B (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__A_N (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__B (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__C_N (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__B (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__A (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__A_N (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__B (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__C_N (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A2 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__A2 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A2 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__B1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__B1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__B (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__B1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__B (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__B1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__B1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__B1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__B1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__B1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A2 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__A2 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__B1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__B1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__B1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A2 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A2 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__A2 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A2 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__C (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A3 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A3 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__A3 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__A2 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__C (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__A3 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A3 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__B (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__B (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A2 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__B (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__B (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A0 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A1 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__C1 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__A3 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A2 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A1 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__B (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A3 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A0 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__B (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__B (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A3 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A3 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__B1 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A2 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A2 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A3 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__B (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A1 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A2 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__B (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__B (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A2 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A3 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A1 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__S0 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__A (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__A (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__S (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__S0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__S0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__A (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6237__A (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A1 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__B1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__B1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__B1 (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__B (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A3 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__B (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A2 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A0 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A2 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A0 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__B2 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__B2 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A2 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A2 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A3 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__B1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A2 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__B1 (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__B1 (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A3 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__B1 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A2 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A2 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__B1 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__B1 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__B2 (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__B2 (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A3 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__B1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__B (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A2 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__B (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__A2 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A2 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__B2 (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__B2 (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__C (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__B1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A0 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A2 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A2 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__B (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__B (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__B1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__B1 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__B (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__B (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__B (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__B2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__B2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__B1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__B1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__B2 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__B2 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__C (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__B (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__B (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A3 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A2 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__B (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__B (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__B1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__B (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__B1 (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A4 (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__C1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__B (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A3 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A0 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A1_N (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__B (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A2 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__B (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__B (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__B (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A0 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__A1 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__B (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__B (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A1 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__B (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__B1 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__B (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__C (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__B (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__B1 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__A2 (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__A2 (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A2 (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A2 (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__B2 (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A3 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A3 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__D (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__A (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__B1 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__B (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A3 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__C (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__B1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A0 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__B (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__B (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__A0 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__B1 (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__B (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__C (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A2 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__A1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__B (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A2 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A2 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__B (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__B (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__B (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A0 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__B (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A3 (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A2 (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__B (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A2 (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__B (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__B (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A2 (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A1 (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A1 (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__C (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__A (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__A (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__A (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__B (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__B (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__C1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__C1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__C1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__C1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__B2 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__B2 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__A2 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A2 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A2 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A2 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A2 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A2 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A2 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A2 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A2 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A2 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A1 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__A (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A2 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__C (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A2 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A2 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A1 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__B1 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A2 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A1 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__B (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__C1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__B1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__C (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__C_N (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__A3 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A2 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__A (.DIODE(_1715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__B (.DIODE(_1715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__C (.DIODE(_1715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__B1 (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__B1 (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__B1 (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__B1 (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__B1 (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__B (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__B (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__D (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A1 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A1 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__B (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__C1 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A2 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__S (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A1 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__S (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__S (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__S (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__S (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__B (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A2 (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__S (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__S (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A3 (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A2 (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A2 (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__C (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A2 (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A2 (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__C (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__C (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__C (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__C (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__C (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__C (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__B (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__B1 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A1 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__S (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__A (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A1 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A1 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A1 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__B1 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A1 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A1 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__D1 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A2 (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A0 (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A2 (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__B (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__B (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__B (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A0 (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A0 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A2 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__B (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__B (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A0 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A1 (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A2 (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__B (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A2 (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A1 (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__B2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__B1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__A2 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__C1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A2 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__B2 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__B1 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__A3 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A0 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A0 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__B (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__B (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A0 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__B (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__B (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__A2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A2 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__B (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B2 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__B1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__A (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__B1 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__S0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__S (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A1 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__B (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__B (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__S0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__S (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A2 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A2 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__B1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__A2 (.DIODE(_1767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__B1 (.DIODE(_1767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__A2 (.DIODE(_1767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__B (.DIODE(_1767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A1 (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__B1 (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__B2 (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__B1 (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__C (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__B1 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A1 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A1 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A1 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__B1 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__D (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A2 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__B2 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__B2 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__B2 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__B2 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A2 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__B2 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__B2 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__B (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__B (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__B (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__S (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A0 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A0 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__S (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__S (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__S (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__S (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__C1 (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__B (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A1 (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__B (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__A (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__A (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__S (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__S (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__S (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__A2 (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__A2 (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A2 (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__B1 (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__B2 (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__B2 (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__S (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__B2 (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__B2 (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__C1 (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__B2 (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__C1 (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__C1 (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__C1 (.DIODE(_1795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A2 (.DIODE(_1795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__A2 (.DIODE(_1795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__B (.DIODE(_1795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__A2 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A2 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__C (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A2 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A1 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__A (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__C (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A1 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__B (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__A (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__B (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A1 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A1 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A1 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__A (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A1 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__A (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__A (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__S (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__C1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__S (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__A1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__C1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A2 (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A2 (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__A2 (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A2 (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A2 (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A2 (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A2 (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__B (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__B (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__B (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__C1 (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__C1 (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__C1 (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__C1 (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__C1 (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__C1 (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__C1 (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__C1 (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__C1 (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__C1 (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__A (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__S (.DIODE(_1835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__S (.DIODE(_1835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__S (.DIODE(_1835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A (.DIODE(_1835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A (.DIODE(_1835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A (.DIODE(_1835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A (.DIODE(_1835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A (.DIODE(_1835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__B (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__C1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__B1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__C1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__S (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__S (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__S (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__S (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__S (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A2 (.DIODE(_1838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A (.DIODE(_1838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A (.DIODE(_1838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A (.DIODE(_1838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A2 (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A2 (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A1 (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A1 (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__B2 (.DIODE(_1841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A3 (.DIODE(_1841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__B1 (.DIODE(_1841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A1 (.DIODE(_1841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A2 (.DIODE(_1841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A2 (.DIODE(_1841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__B (.DIODE(_1841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A1 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A2 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__A (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__B1 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__C (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__B1 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A2 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__B (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__C (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A1 (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A_N (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__C (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__B1 (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A2 (.DIODE(_1886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A2 (.DIODE(_1886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A2 (.DIODE(_1886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A2 (.DIODE(_1886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__S (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A1 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__B1 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B1 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A0 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__B (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A2 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A2 (.DIODE(_1902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__B2 (.DIODE(_1902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A1 (.DIODE(_1902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__A2 (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__B1 (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__B1 (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__B (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A3 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__B (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__A1 (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A2 (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__B1 (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__C (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__B1 (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A2 (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A0 (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__B (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__S (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__S (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__S (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A1 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__S (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__S (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__S0 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__S0 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__S (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__B (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__B (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__B (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__B1 (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A1 (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__S1 (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1_N (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__S1 (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__B2 (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A1 (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__B (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__S (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__B (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__B (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__A (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__S (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__S (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__S0 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__B2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__S (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__A0 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__B (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__B (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__B1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__B (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B (.DIODE(_2018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__B (.DIODE(_2018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A0 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__C (.DIODE(_2027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__B (.DIODE(_2027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__B (.DIODE(_2027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A0 (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__D (.DIODE(_2033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__B (.DIODE(_2033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__C (.DIODE(_2033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__B1 (.DIODE(_2033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A0 (.DIODE(_2036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__S (.DIODE(_2044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__S (.DIODE(_2044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__S (.DIODE(_2044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__S (.DIODE(_2044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__S (.DIODE(_2044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__S (.DIODE(_2044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__S (.DIODE(_2044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__S (.DIODE(_2044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__S (.DIODE(_2044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__S (.DIODE(_2044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__C (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__C (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__C (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__C (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__C (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__B (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__B1 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__B1 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__B1 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B1 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__B1 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__B1 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A2 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__B1 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__B (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__B1 (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__B1 (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B1 (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__B1 (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__B (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__S (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__B1 (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__B1 (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__B1 (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__B1 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A1 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__S (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__B1 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A1 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__S (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A1 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__S (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__S (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__S (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__S (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__S (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__S (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__S (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__S (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__S (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__S (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__S (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__S (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__S (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__C (.DIODE(_2099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__B (.DIODE(_2099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A3 (.DIODE(_2102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__B2 (.DIODE(_2102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A4 (.DIODE(_2102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__C (.DIODE(_2102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__B1 (.DIODE(_2102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__B1 (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A2_N (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__B2 (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A2 (.DIODE(_2126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B1 (.DIODE(_2126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A2 (.DIODE(_2128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__B1 (.DIODE(_2128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A2 (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__A (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__B1 (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__B1 (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__B1 (.DIODE(_2133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__B (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__B (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A2 (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A1 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A1 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A1 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A1 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__A1 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A1 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A1 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B2 (.DIODE(_2137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A0 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A0 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__B2 (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__B2 (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__B2 (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__B2 (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__B2 (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__B2 (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__B2 (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__B2 (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__B2 (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A1 (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A1 (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__B1 (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A1 (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A1 (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A1 (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B1 (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A1 (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__C1 (.DIODE(_2183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A (.DIODE(_2184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A (.DIODE(_2184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__B (.DIODE(_2184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__B2 (.DIODE(_2186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A2 (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A0 (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A2 (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__B1 (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__B1 (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__B1 (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B1 (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__B1 (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__B1 (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B1 (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__B1 (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__B1 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A1 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__B1 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A2 (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A2 (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__B (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__A (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__A3 (.DIODE(_2231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B1 (.DIODE(_2231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__C (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__B (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__B2 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A2 (.DIODE(_2241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A0 (.DIODE(_2241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B2 (.DIODE(_2241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__D (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A (.DIODE(_2263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A_N (.DIODE(_2263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A2 (.DIODE(_2263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__B (.DIODE(_2266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A0 (.DIODE(_2266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A2 (.DIODE(_2266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A2 (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__B (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A2 (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__B (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__B (.DIODE(_2295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A (.DIODE(_2295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A2 (.DIODE(_2295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__B2 (.DIODE(_2297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__A2 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A0 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A0 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__B1_N (.DIODE(_2303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__C_N (.DIODE(_2303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A2 (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A2 (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__A2 (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A2 (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A2 (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A2 (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A2 (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A2 (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A2 (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A2 (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A2 (.DIODE(_2315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__B (.DIODE(_2315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__B (.DIODE(_2315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__A2 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A0 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__B (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__S (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__S (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__S (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__S (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__S (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__S (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__S (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__S (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__S (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__S (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__B2 (.DIODE(_2356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__B (.DIODE(_2364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A (.DIODE(_2364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A2 (.DIODE(_2364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__A2 (.DIODE(_2367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A0 (.DIODE(_2367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A2 (.DIODE(_2367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__B (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A2 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A2 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A2 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A2 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A2 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A2 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A2 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A2 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__A2 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__C (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__B1 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__B1 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__B1 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__B1 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__B1 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__B1 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__B1 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B1 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__B1 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__B1 (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__B_N (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B1 (.DIODE(_2394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__A2 (.DIODE(_2396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A0 (.DIODE(_2396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A0 (.DIODE(_2396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__B1 (.DIODE(_2415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A1 (.DIODE(_2419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__B (.DIODE(_2419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A1 (.DIODE(_2419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__B1 (.DIODE(_2425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__A2 (.DIODE(_2427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A0 (.DIODE(_2427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__B (.DIODE(_2427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__B1 (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__B1 (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__C1 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A2 (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__B (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A0 (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A2 (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__B1 (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__B1 (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__C1 (.DIODE(_2499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__B1_N (.DIODE(_2499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__B1 (.DIODE(_2513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__B1 (.DIODE(_2523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A0 (.DIODE(_2523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__B (.DIODE(_2523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__C1 (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__C1 (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__C1 (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__B (.DIODE(_2539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A2 (.DIODE(_2539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__B (.DIODE(_2539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__C1 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A2 (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__B (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A2 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__B2 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__B1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A1 (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__A2 (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A0 (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A0 (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__B (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A2 (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A0 (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__B (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__A2 (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__A2 (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A0 (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A2 (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A2 (.DIODE(_2620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__B (.DIODE(_2620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__S (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__S (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__S (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__S (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__S (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__S (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__S (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__S (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__S (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__S (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__S (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__S (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__S (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__S (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__S (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__S (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__S (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__S (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__S (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__S (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__B (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__B (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__B (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__B (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__B (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__B (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A1 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A1 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A1 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A1 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A1 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A1 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A1 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A1 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A2 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__B (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__B (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__B (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__B (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__C1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__C1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__C1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__C1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__C1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__C1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__C1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__C1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__C1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__C1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A2 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__A1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__A1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__A1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__A1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A2 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A2 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__A1 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A1 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A1 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A1 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A1 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A1 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A1 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A2 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A1 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A1 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A1 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__A1 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__A1 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A1 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A1 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A2 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__A1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__A1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A2 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A2 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__B (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__A (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__A (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__A (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__A (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__B (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__B (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__A (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__A (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__A (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__A (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__B (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__A (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__B (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__A (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__A (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__B (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__A (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__A (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__A (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__A (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__B (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__B (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__B (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__B (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__B (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__C1 (.DIODE(_2726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__C1 (.DIODE(_2726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__C1 (.DIODE(_2726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__C1 (.DIODE(_2726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__C1 (.DIODE(_2726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__C1 (.DIODE(_2726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__C1 (.DIODE(_2726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__C1 (.DIODE(_2726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__C1 (.DIODE(_2726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__C1 (.DIODE(_2726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__C1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__C1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__C1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__C1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__C1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__C1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__C1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__C1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__C1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__C1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A2 (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A2 (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A2 (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A2 (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A2 (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__A2 (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A2 (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A2 (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__A (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__B (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__B (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__B (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__B (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__A (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A2 (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A2 (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A2 (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A2 (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A2 (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A2 (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__A2 (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__B (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A2 (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__B (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__C1 (.DIODE(_2753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__C1 (.DIODE(_2753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__C1 (.DIODE(_2753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__C1 (.DIODE(_2753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__C1 (.DIODE(_2753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__C1 (.DIODE(_2753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__C1 (.DIODE(_2753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__C1 (.DIODE(_2753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__C1 (.DIODE(_2753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__C1 (.DIODE(_2753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__A2 (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A2 (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__A2 (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A2 (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A2 (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__A2 (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A2 (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A2 (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__B (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__B (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__B (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__B (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__B (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__B (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__B (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__B (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__B (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__B (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__B (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__B (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__B (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__B (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__C1 (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__C1 (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__C1 (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__C1 (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__C1 (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__C1 (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__C1 (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__C1 (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__C1 (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__C1 (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__C1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__C1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__C1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__C1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__C1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__C1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__C1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__C1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__C1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__C1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A2 (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A2 (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__A2 (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A2 (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A2 (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__A2 (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A2 (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__A2 (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__B (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__B (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__B (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__B (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__C1 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__C1 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__C1 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__C1 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__C1 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__C1 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__C1 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__C1 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__C1 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__C1 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__A2 (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__A2 (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A2 (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A2 (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__A2 (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A2 (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A2 (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A2 (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__A (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__B (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__B (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__B (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__B (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__C1 (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__C1 (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__C1 (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__C1 (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__C1 (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__C1 (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__C1 (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__C1 (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__C1 (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__C1 (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__C1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__C1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__C1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__C1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__C1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__C1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__C1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__C1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__C1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__C1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A2 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__A2 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A2 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A2 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A2 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A2 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A2 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__A2 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__C1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__C1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__C1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__C1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__C1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__C1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__C1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__C1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__C1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__C1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__A2 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A2 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A2 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A2 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A2 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A2 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A2 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__B (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A2 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__B (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__C1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__C1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__C1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__C1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__C1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__C1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__C1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__C1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__C1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__C1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__B (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__B (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__B (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__B (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__A (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__C1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__C1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__C1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__C1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__C1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__C1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__C1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__C1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__C1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__C1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__B1 (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__B1 (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__B1 (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__B1 (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__C1 (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__C1 (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__A (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__A (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__B1 (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__B1 (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__A (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A1 (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A1 (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A1 (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__A (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__A1 (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__B1 (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__A1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__A1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__B1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__A1 (.DIODE(_2892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__A1 (.DIODE(_2892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__A1 (.DIODE(_2892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__B2 (.DIODE(_2892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A1 (.DIODE(_2892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__B2 (.DIODE(_2892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A1 (.DIODE(_2892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__B1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__B1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__B1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__B1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__B1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A2 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__S (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__B1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__A2 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__B1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__A2 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A2 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A2 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A2 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A2 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A2 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A2 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__B (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__A2 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A2 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A3 (.DIODE(_2901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__B1 (.DIODE(_2901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A0 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__B (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__C (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A2 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__S (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__A2 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A2 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__S (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A2 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__S (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A2 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A1 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__B (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__B (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__B (.DIODE(_2992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__B (.DIODE(_2992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__B (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__B (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__B (.DIODE(_3027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__B (.DIODE(_3027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A3 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A3 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__C (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A3 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__A3 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A3 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__A3 (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A3 (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__A3 (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__C (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A3 (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__A3 (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__A3 (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__B2 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__A (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__A (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__B2 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__B2 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__B2 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__A2 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__A2 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__B2 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__B2 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A2 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__B2 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__B2 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__A (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__A (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__A (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__A (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__A (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__C (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A1 (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__B_N (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__A2_N (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__A2_N (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A2_N (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__A2_N (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__A2_N (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A2_N (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__A2_N (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__C (.DIODE(_3105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__C (.DIODE(_3117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A2 (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__C (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__B (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__B (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__B1 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__B1 (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__B1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A1 (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__B (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__B (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__B1 (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__S (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__S (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__B (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__C (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__A2 (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__C1 (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__B (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__C1 (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__B (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__S (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__A2 (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__A2 (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__A3 (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__S (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__S (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__S (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__S (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__S (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__S (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A2 (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__S (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__S (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__S (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__S (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__S (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__S (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__S (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__S (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__S (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__S (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__S (.DIODE(_3231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__S (.DIODE(_3231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__S (.DIODE(_3231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__S (.DIODE(_3231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__S (.DIODE(_3231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__S (.DIODE(_3231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__A (.DIODE(_3231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__S (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__S (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__S (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__S (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__S (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__S (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__S (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__S (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__S (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__S (.DIODE(_3232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__A (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__A (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__A (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A0 (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__A (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__A (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__A (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__A (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A0 (.DIODE(_3289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A2 (.DIODE(_3298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A2 (.DIODE(_3298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A2 (.DIODE(_3298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__B (.DIODE(_3298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__B (.DIODE(_3310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A2 (.DIODE(_3310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__B (.DIODE(_3310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__B (.DIODE(_3310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__B (.DIODE(_3310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__B (.DIODE(_3310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A2 (.DIODE(_3310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A2 (.DIODE(_3310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__A2 (.DIODE(_3310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A (.DIODE(_3310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__A2 (.DIODE(_3311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A2 (.DIODE(_3311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A2 (.DIODE(_3311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A2 (.DIODE(_3311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A2 (.DIODE(_3311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A2 (.DIODE(_3311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__A2 (.DIODE(_3311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__A2 (.DIODE(_3311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__A2 (.DIODE(_3311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A2 (.DIODE(_3311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__C1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__C1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__C1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__C1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__C1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__C1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__C1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__C1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__C1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__C1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__C1 (.DIODE(_3332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__C1 (.DIODE(_3332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__C1 (.DIODE(_3332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__C1 (.DIODE(_3332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__C1 (.DIODE(_3332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__C1 (.DIODE(_3332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__C1 (.DIODE(_3332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__C1 (.DIODE(_3332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__C1 (.DIODE(_3332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__C1 (.DIODE(_3332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__S (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__A2 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__B1 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__A2 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__A (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__S (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__S (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__S (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__B1 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__B (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__S (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__S (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A2 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__C1 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__S (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__S (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__S (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__S (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A2 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__S (.DIODE(_3387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A (.DIODE(_3387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__A (.DIODE(_3387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__A (.DIODE(_3387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__A (.DIODE(_3387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A (.DIODE(_3387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__S (.DIODE(_3390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__S (.DIODE(_3390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__S (.DIODE(_3390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__S (.DIODE(_3390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__S (.DIODE(_3390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__S (.DIODE(_3390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__S (.DIODE(_3390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__S (.DIODE(_3390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A0 (.DIODE(\core_0.de_jmp_pred ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A (.DIODE(\core_0.de_jmp_pred ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A2 (.DIODE(\core_0.de_jmp_pred ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__B2 (.DIODE(\core_0.dec_jump_cond_code[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A1 (.DIODE(\core_0.dec_jump_cond_code[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__D (.DIODE(\core_0.dec_jump_cond_code[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__A (.DIODE(\core_0.dec_jump_cond_code[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__A2 (.DIODE(\core_0.dec_jump_cond_code[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__B (.DIODE(\core_0.dec_jump_cond_code[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__B2 (.DIODE(\core_0.dec_jump_cond_code[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A1 (.DIODE(\core_0.dec_jump_cond_code[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A2 (.DIODE(\core_0.dec_jump_cond_code[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__C (.DIODE(\core_0.dec_jump_cond_code[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__S (.DIODE(\core_0.dec_jump_cond_code[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A2 (.DIODE(\core_0.dec_jump_cond_code[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__C (.DIODE(\core_0.dec_jump_cond_code[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A (.DIODE(\core_0.dec_jump_cond_code[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__B2 (.DIODE(\core_0.dec_jump_cond_code[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__B1 (.DIODE(\core_0.dec_jump_cond_code[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__B (.DIODE(\core_0.dec_jump_cond_code[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__B1 (.DIODE(\core_0.dec_jump_cond_code[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__C1 (.DIODE(\core_0.dec_jump_cond_code[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__B2 (.DIODE(\core_0.dec_jump_cond_code[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__S (.DIODE(\core_0.dec_jump_cond_code[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__A1 (.DIODE(\core_0.dec_jump_cond_code[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__A1 (.DIODE(\core_0.dec_jump_cond_code[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__A1 (.DIODE(\core_0.dec_jump_cond_code[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__B2 (.DIODE(\core_0.dec_jump_cond_code[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__C_N (.DIODE(\core_0.dec_jump_cond_code[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A1 (.DIODE(\core_0.dec_jump_cond_code[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A1 (.DIODE(\core_0.dec_jump_cond_code[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__B (.DIODE(\core_0.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__B (.DIODE(\core_0.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__D (.DIODE(\core_0.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A_N (.DIODE(\core_0.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__C (.DIODE(\core_0.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__B (.DIODE(\core_0.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A_N (.DIODE(\core_0.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__A (.DIODE(\core_0.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A (.DIODE(\core_0.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A (.DIODE(\core_0.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A0 (.DIODE(\core_0.dec_mem_we ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A1 (.DIODE(\core_0.dec_mem_we ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__A2 (.DIODE(\core_0.dec_pc_inc ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__B1 (.DIODE(\core_0.dec_pc_inc ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A1 (.DIODE(\core_0.dec_pc_inc ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__B (.DIODE(\core_0.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A1 (.DIODE(\core_0.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__B (.DIODE(\core_0.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__B (.DIODE(\core_0.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A1 (.DIODE(\core_0.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(\core_0.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__B (.DIODE(\core_0.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A (.DIODE(\core_0.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__A (.DIODE(\core_0.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__A2 (.DIODE(\core_0.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__C1 (.DIODE(\core_0.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A (.DIODE(\core_0.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A (.DIODE(\core_0.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__D1 (.DIODE(\core_0.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A (.DIODE(\core_0.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A (.DIODE(\core_0.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A (.DIODE(\core_0.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__B1 (.DIODE(\core_0.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__B2 (.DIODE(\core_0.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__A (.DIODE(\core_0.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A (.DIODE(\core_0.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__A (.DIODE(\core_0.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A (.DIODE(\core_0.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__B (.DIODE(\core_0.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A (.DIODE(\core_0.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A1 (.DIODE(\core_0.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A1 (.DIODE(\core_0.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A1 (.DIODE(\core_0.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__B (.DIODE(\core_0.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A1 (.DIODE(\core_0.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__B (.DIODE(\core_0.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__B (.DIODE(\core_0.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A (.DIODE(\core_0.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__B (.DIODE(\core_0.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__B (.DIODE(\core_0.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__A1 (.DIODE(\core_0.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A1 (.DIODE(\core_0.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A1 (.DIODE(\core_0.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__B2 (.DIODE(\core_0.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A1 (.DIODE(\core_0.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__B2 (.DIODE(\core_0.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A1 (.DIODE(\core_0.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A1 (.DIODE(\core_0.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__B2 (.DIODE(\core_0.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A1 (.DIODE(\core_0.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A1 (.DIODE(\core_0.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__B2 (.DIODE(\core_0.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__A1 (.DIODE(\core_0.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A1 (.DIODE(\core_0.decode.i_instr_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__B (.DIODE(\core_0.decode.i_instr_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__B (.DIODE(\core_0.decode.i_instr_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__B (.DIODE(\core_0.decode.i_instr_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__B (.DIODE(\core_0.decode.i_instr_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__B_N (.DIODE(\core_0.decode.i_instr_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A_N (.DIODE(\core_0.decode.i_instr_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A1 (.DIODE(\core_0.decode.i_instr_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A (.DIODE(\core_0.decode.i_instr_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A (.DIODE(\core_0.decode.i_instr_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A (.DIODE(\core_0.decode.i_instr_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__A (.DIODE(\core_0.decode.i_instr_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A (.DIODE(\core_0.decode.i_instr_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__B (.DIODE(\core_0.decode.i_instr_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A (.DIODE(\core_0.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A (.DIODE(\core_0.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A1 (.DIODE(\core_0.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A (.DIODE(\core_0.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A (.DIODE(\core_0.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__B (.DIODE(\core_0.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A1 (.DIODE(\core_0.decode.oc_alu_mode[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__B1 (.DIODE(\core_0.decode.oc_alu_mode[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A1 (.DIODE(\core_0.decode.oc_alu_mode[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A1 (.DIODE(\core_0.decode.oc_alu_mode[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__A (.DIODE(\core_0.decode.oc_alu_mode[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A2 (.DIODE(\core_0.decode.oc_alu_mode[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A (.DIODE(\core_0.decode.oc_alu_mode[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A (.DIODE(\core_0.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__D (.DIODE(\core_0.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__B (.DIODE(\core_0.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__C1 (.DIODE(\core_0.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__B1 (.DIODE(\core_0.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__A (.DIODE(\core_0.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A1 (.DIODE(\core_0.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A (.DIODE(\core_0.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A (.DIODE(\core_0.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A1 (.DIODE(\core_0.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A1 (.DIODE(\core_0.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A1 (.DIODE(\core_0.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A1 (.DIODE(\core_0.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__B2 (.DIODE(\core_0.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A1 (.DIODE(\core_0.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__A1 (.DIODE(\core_0.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__D (.DIODE(\core_0.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A (.DIODE(\core_0.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A (.DIODE(\core_0.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A (.DIODE(\core_0.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A (.DIODE(\core_0.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__C (.DIODE(\core_0.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A1 (.DIODE(\core_0.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A (.DIODE(\core_0.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__B2 (.DIODE(\core_0.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__A (.DIODE(\core_0.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A1 (.DIODE(\core_0.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A (.DIODE(\core_0.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__B2 (.DIODE(\core_0.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B2 (.DIODE(\core_0.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A (.DIODE(\core_0.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__C1 (.DIODE(\core_0.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__B2 (.DIODE(\core_0.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__B2 (.DIODE(\core_0.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__B (.DIODE(\core_0.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A (.DIODE(\core_0.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__B1 (.DIODE(\core_0.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A1 (.DIODE(\core_0.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A1 (.DIODE(\core_0.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A1 (.DIODE(\core_0.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__B1 (.DIODE(\core_0.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A1 (.DIODE(\core_0.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A1 (.DIODE(\core_0.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__C (.DIODE(\core_0.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A (.DIODE(\core_0.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__B2 (.DIODE(\core_0.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__C1 (.DIODE(\core_0.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__B2 (.DIODE(\core_0.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__C1 (.DIODE(\core_0.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A1 (.DIODE(\core_0.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__B2 (.DIODE(\core_0.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__A1 (.DIODE(\core_0.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A (.DIODE(\core_0.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A (.DIODE(\core_0.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__A0 (.DIODE(\core_0.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(\core_0.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A0 (.DIODE(\core_0.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A (.DIODE(\core_0.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A (.DIODE(\core_0.ew_data[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1 (.DIODE(\core_0.ew_data[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A1 (.DIODE(\core_0.ew_data[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A (.DIODE(\core_0.ew_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A1 (.DIODE(\core_0.ew_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A1 (.DIODE(\core_0.ew_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A0 (.DIODE(\core_0.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A1 (.DIODE(\core_0.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__A0 (.DIODE(\core_0.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A (.DIODE(\core_0.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A0 (.DIODE(\core_0.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A1 (.DIODE(\core_0.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A0 (.DIODE(\core_0.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__A (.DIODE(\core_0.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A0 (.DIODE(\core_0.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__A1 (.DIODE(\core_0.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A0 (.DIODE(\core_0.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A (.DIODE(\core_0.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A0 (.DIODE(\core_0.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A1 (.DIODE(\core_0.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A0 (.DIODE(\core_0.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A (.DIODE(\core_0.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A0 (.DIODE(\core_0.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A1 (.DIODE(\core_0.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A0 (.DIODE(\core_0.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A (.DIODE(\core_0.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A0 (.DIODE(\core_0.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__A1 (.DIODE(\core_0.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A0 (.DIODE(\core_0.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A (.DIODE(\core_0.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A0 (.DIODE(\core_0.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A1 (.DIODE(\core_0.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A0 (.DIODE(\core_0.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A (.DIODE(\core_0.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A (.DIODE(\core_0.ew_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A1 (.DIODE(\core_0.ew_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A1 (.DIODE(\core_0.ew_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A_N (.DIODE(\core_0.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1 (.DIODE(\core_0.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__B_N (.DIODE(\core_0.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__B (.DIODE(\core_0.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A (.DIODE(\core_0.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A (.DIODE(\core_0.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A1 (.DIODE(\core_0.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A2 (.DIODE(\core_0.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A1 (.DIODE(\core_0.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__B (.DIODE(\core_0.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A (.DIODE(\core_0.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A (.DIODE(\core_0.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A1 (.DIODE(\core_0.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A3 (.DIODE(\core_0.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__B2 (.DIODE(\core_0.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A3 (.DIODE(\core_0.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A (.DIODE(\core_0.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A (.DIODE(\core_0.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A1 (.DIODE(\core_0.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A0 (.DIODE(\core_0.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A0 (.DIODE(\core_0.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A3 (.DIODE(\core_0.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A (.DIODE(\core_0.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A (.DIODE(\core_0.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A1 (.DIODE(\core_0.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A1 (.DIODE(\core_0.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A1 (.DIODE(\core_0.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A0 (.DIODE(\core_0.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__A (.DIODE(\core_0.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A (.DIODE(\core_0.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A1 (.DIODE(\core_0.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A3 (.DIODE(\core_0.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__B2 (.DIODE(\core_0.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A2 (.DIODE(\core_0.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A0 (.DIODE(\core_0.ew_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__S (.DIODE(\core_0.ew_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__B2 (.DIODE(\core_0.ew_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A1 (.DIODE(\core_0.ew_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__A1 (.DIODE(\core_0.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A (.DIODE(\core_0.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__B (.DIODE(\core_0.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A1 (.DIODE(\core_0.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__B (.DIODE(\core_0.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A (.DIODE(\core_0.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__A1 (.DIODE(\core_0.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__B2 (.DIODE(\core_0.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A (.DIODE(\core_0.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A (.DIODE(\core_0.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__B1 (.DIODE(\core_0.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A0 (.DIODE(\core_0.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A0 (.DIODE(\core_0.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B2 (.DIODE(\core_0.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A1 (.DIODE(\core_0.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A (.DIODE(\core_0.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A (.DIODE(\core_0.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A (.DIODE(\core_0.execute.alu_flag_reg.o_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__B2 (.DIODE(\core_0.execute.alu_flag_reg.o_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A (.DIODE(\core_0.execute.alu_flag_reg.o_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A (.DIODE(\core_0.execute.alu_flag_reg.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__B2 (.DIODE(\core_0.execute.alu_flag_reg.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A1 (.DIODE(\core_0.execute.alu_flag_reg.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__B1 (.DIODE(\core_0.execute.alu_mul_div.comp ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A (.DIODE(\core_0.execute.alu_mul_div.comp ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A (.DIODE(\core_0.execute.alu_mul_div.comp ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A (.DIODE(\core_0.execute.alu_mul_div.comp ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A2 (.DIODE(\core_0.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A0 (.DIODE(\core_0.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__B1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__A1_N (.DIODE(\core_0.execute.alu_mul_div.div_cur[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__A0 (.DIODE(\core_0.execute.alu_mul_div.div_cur[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A0 (.DIODE(\core_0.execute.alu_mul_div.div_cur[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A0 (.DIODE(\core_0.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__A0 (.DIODE(\core_0.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A0 (.DIODE(\core_0.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A0 (.DIODE(\core_0.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A1 (.DIODE(\core_0.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__A (.DIODE(\core_0.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__B1 (.DIODE(\core_0.execute.alu_mul_div.div_res[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A1 (.DIODE(\core_0.execute.alu_mul_div.div_res[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__B1 (.DIODE(\core_0.execute.alu_mul_div.div_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A1 (.DIODE(\core_0.execute.alu_mul_div.div_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__B1 (.DIODE(\core_0.execute.alu_mul_div.div_res[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A1 (.DIODE(\core_0.execute.alu_mul_div.div_res[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__B1 (.DIODE(\core_0.execute.alu_mul_div.div_res[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A1 (.DIODE(\core_0.execute.alu_mul_div.div_res[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__B1 (.DIODE(\core_0.execute.alu_mul_div.div_res[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A1 (.DIODE(\core_0.execute.alu_mul_div.div_res[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__B1 (.DIODE(\core_0.execute.alu_mul_div.div_res[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A1 (.DIODE(\core_0.execute.alu_mul_div.div_res[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__B1 (.DIODE(\core_0.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__A2_N (.DIODE(\core_0.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A2 (.DIODE(\core_0.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A2 (.DIODE(\core_0.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A2 (.DIODE(\core_0.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A2 (.DIODE(\core_0.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__C1 (.DIODE(\core_0.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A (.DIODE(\core_0.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A (.DIODE(\core_0.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__B (.DIODE(\core_0.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A1 (.DIODE(\core_0.execute.alu_mul_div.mul_res[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A (.DIODE(\core_0.execute.alu_mul_div.mul_res[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__A (.DIODE(\core_0.execute.alu_mul_div.mul_res[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A2 (.DIODE(\core_0.execute.alu_mul_div.mul_res[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__B2 (.DIODE(\core_0.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__A (.DIODE(\core_0.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A (.DIODE(\core_0.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A2 (.DIODE(\core_0.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__A1 (.DIODE(\core_0.execute.alu_mul_div.mul_res[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A (.DIODE(\core_0.execute.alu_mul_div.mul_res[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__A (.DIODE(\core_0.execute.alu_mul_div.mul_res[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A2 (.DIODE(\core_0.execute.alu_mul_div.mul_res[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__A0 (.DIODE(\core_0.execute.alu_mul_div.mul_res[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A (.DIODE(\core_0.execute.alu_mul_div.mul_res[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A2 (.DIODE(\core_0.execute.alu_mul_div.mul_res[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A1 (.DIODE(\core_0.execute.alu_mul_div.mul_res[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A (.DIODE(\core_0.execute.alu_mul_div.mul_res[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__A (.DIODE(\core_0.execute.alu_mul_div.mul_res[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A0 (.DIODE(\core_0.execute.alu_mul_div.mul_res[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A1 (.DIODE(\core_0.execute.alu_mul_div.mul_res[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A_N (.DIODE(\core_0.execute.alu_mul_div.mul_res[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__B (.DIODE(\core_0.execute.alu_mul_div.mul_res[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A2 (.DIODE(\core_0.execute.alu_mul_div.mul_res[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A0 (.DIODE(\core_0.execute.alu_mul_div.mul_res[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A (.DIODE(\core_0.execute.alu_mul_div.mul_res[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A2 (.DIODE(\core_0.execute.alu_mul_div.mul_res[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__A1 (.DIODE(\core_0.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A1 (.DIODE(\core_0.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__B1 (.DIODE(\core_0.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A1 (.DIODE(\core_0.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__B1 (.DIODE(\core_0.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__A1 (.DIODE(\core_0.execute.pc_high_buff_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__A0 (.DIODE(\core_0.execute.pc_high_buff_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A1 (.DIODE(\core_0.execute.pc_high_buff_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__A1 (.DIODE(\core_0.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__B1 (.DIODE(\core_0.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A1 (.DIODE(\core_0.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__A1 (.DIODE(\core_0.execute.pc_high_buff_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__A1 (.DIODE(\core_0.execute.pc_high_buff_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A1 (.DIODE(\core_0.execute.pc_high_buff_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A1 (.DIODE(\core_0.execute.pc_high_buff_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__A1 (.DIODE(\core_0.execute.pc_high_buff_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A1 (.DIODE(\core_0.execute.pc_high_buff_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__A1 (.DIODE(\core_0.execute.pc_high_buff_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__A1 (.DIODE(\core_0.execute.pc_high_buff_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A1 (.DIODE(\core_0.execute.pc_high_buff_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__A (.DIODE(\core_0.execute.pc_high_buff_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__A0 (.DIODE(\core_0.execute.pc_high_buff_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A1 (.DIODE(\core_0.execute.pc_high_buff_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__A3 (.DIODE(\core_0.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__D (.DIODE(\core_0.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__A2 (.DIODE(\core_0.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__B (.DIODE(\core_0.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A1 (.DIODE(\core_0.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A (.DIODE(\core_0.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(\core_0.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__A (.DIODE(\core_0.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__A2 (.DIODE(\core_0.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__C (.DIODE(\core_0.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__A0 (.DIODE(\core_0.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__A1 (.DIODE(\core_0.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__A (.DIODE(\core_0.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A (.DIODE(\core_0.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__A (.DIODE(\core_0.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__A0 (.DIODE(\core_0.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__B1 (.DIODE(\core_0.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A (.DIODE(\core_0.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A1 (.DIODE(\core_0.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A (.DIODE(\core_0.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__A1 (.DIODE(\core_0.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__B (.DIODE(\core_0.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__A1 (.DIODE(\core_0.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__A1 (.DIODE(\core_0.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A1 (.DIODE(\core_0.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__B2 (.DIODE(\core_0.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A (.DIODE(\core_0.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A (.DIODE(\core_0.execute.rf.reg_outputs[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__C_N (.DIODE(\core_0.execute.rf.reg_outputs[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__D (.DIODE(\core_0.execute.rf.reg_outputs[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A (.DIODE(\core_0.execute.rf.reg_outputs[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__A (.DIODE(\core_0.execute.rf.reg_outputs[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__B2 (.DIODE(\core_0.execute.rf.reg_outputs[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A (.DIODE(\core_0.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A1 (.DIODE(\core_0.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A1 (.DIODE(\core_0.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A1 (.DIODE(\core_0.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A (.DIODE(\core_0.execute.rf.reg_outputs[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A1 (.DIODE(\core_0.execute.rf.reg_outputs[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__B2 (.DIODE(\core_0.execute.rf.reg_outputs[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__B2 (.DIODE(\core_0.execute.rf.reg_outputs[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__A (.DIODE(\core_0.execute.rf.reg_outputs[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A1 (.DIODE(\core_0.execute.rf.reg_outputs[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A1 (.DIODE(\core_0.execute.rf.reg_outputs[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__D (.DIODE(\core_0.execute.rf.reg_outputs[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A1 (.DIODE(\core_0.execute.rf.reg_outputs[1][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__A (.DIODE(\core_0.execute.rf.reg_outputs[1][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A1 (.DIODE(\core_0.execute.rf.reg_outputs[1][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A1 (.DIODE(\core_0.execute.rf.reg_outputs[2][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__B2 (.DIODE(\core_0.execute.rf.reg_outputs[2][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__B2 (.DIODE(\core_0.execute.rf.reg_outputs[2][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A1 (.DIODE(\core_0.execute.rf.reg_outputs[2][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__B2 (.DIODE(\core_0.execute.rf.reg_outputs[2][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__A1 (.DIODE(\core_0.execute.rf.reg_outputs[2][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A (.DIODE(\core_0.execute.rf.reg_outputs[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__C (.DIODE(\core_0.execute.rf.reg_outputs[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__D (.DIODE(\core_0.execute.rf.reg_outputs[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__A (.DIODE(\core_0.execute.rf.reg_outputs[3][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__D (.DIODE(\core_0.execute.rf.reg_outputs[3][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__D (.DIODE(\core_0.execute.rf.reg_outputs[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__D (.DIODE(\core_0.execute.rf.reg_outputs[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__D (.DIODE(\core_0.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__A (.DIODE(\core_0.execute.rf.reg_outputs[3][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A (.DIODE(\core_0.execute.rf.reg_outputs[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__C (.DIODE(\core_0.execute.rf.reg_outputs[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__D (.DIODE(\core_0.execute.rf.reg_outputs[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A (.DIODE(\core_0.execute.rf.reg_outputs[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__D (.DIODE(\core_0.execute.rf.reg_outputs[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A (.DIODE(\core_0.execute.rf.reg_outputs[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A (.DIODE(\core_0.execute.rf.reg_outputs[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__D (.DIODE(\core_0.execute.rf.reg_outputs[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__D (.DIODE(\core_0.execute.rf.reg_outputs[3][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__D (.DIODE(\core_0.execute.rf.reg_outputs[3][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__A1 (.DIODE(\core_0.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__D (.DIODE(\core_0.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__A (.DIODE(\core_0.execute.rf.reg_outputs[4][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__C (.DIODE(\core_0.execute.rf.reg_outputs[4][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__B2 (.DIODE(\core_0.execute.rf.reg_outputs[4][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__A (.DIODE(\core_0.execute.rf.reg_outputs[4][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__B2 (.DIODE(\core_0.execute.rf.reg_outputs[4][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A (.DIODE(\core_0.execute.rf.reg_outputs[4][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A (.DIODE(\core_0.execute.rf.reg_outputs[4][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A (.DIODE(\core_0.execute.rf.reg_outputs[4][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__A (.DIODE(\core_0.execute.rf.reg_outputs[4][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__C_N (.DIODE(\core_0.execute.rf.reg_outputs[4][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A (.DIODE(\core_0.execute.rf.reg_outputs[4][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__C (.DIODE(\core_0.execute.rf.reg_outputs[4][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A (.DIODE(\core_0.execute.rf.reg_outputs[4][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A (.DIODE(\core_0.execute.rf.reg_outputs[4][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__B2 (.DIODE(\core_0.execute.rf.reg_outputs[4][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__A (.DIODE(\core_0.execute.rf.reg_outputs[4][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__B2 (.DIODE(\core_0.execute.rf.reg_outputs[4][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A (.DIODE(\core_0.execute.rf.reg_outputs[4][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__B2 (.DIODE(\core_0.execute.rf.reg_outputs[4][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A (.DIODE(\core_0.execute.rf.reg_outputs[4][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A (.DIODE(\core_0.execute.rf.reg_outputs[4][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__C (.DIODE(\core_0.execute.rf.reg_outputs[4][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__B2 (.DIODE(\core_0.execute.rf.reg_outputs[4][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A1 (.DIODE(\core_0.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__B2 (.DIODE(\core_0.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__A (.DIODE(\core_0.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__C (.DIODE(\core_0.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__C (.DIODE(\core_0.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__C (.DIODE(\core_0.execute.rf.reg_outputs[5][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__B2 (.DIODE(\core_0.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__C (.DIODE(\core_0.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__B2 (.DIODE(\core_0.execute.rf.reg_outputs[5][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__B2 (.DIODE(\core_0.execute.rf.reg_outputs[5][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__A (.DIODE(\core_0.execute.rf.reg_outputs[5][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__B2 (.DIODE(\core_0.execute.rf.reg_outputs[5][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A (.DIODE(\core_0.execute.rf.reg_outputs[5][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__B2 (.DIODE(\core_0.execute.rf.reg_outputs[5][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A1 (.DIODE(\core_0.execute.rf.reg_outputs[5][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A (.DIODE(\core_0.execute.rf.reg_outputs[6][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__D (.DIODE(\core_0.execute.rf.reg_outputs[6][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__D (.DIODE(\core_0.execute.rf.reg_outputs[6][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A1 (.DIODE(\core_0.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A1 (.DIODE(\core_0.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__B2 (.DIODE(\core_0.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__A1 (.DIODE(\core_0.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__A1 (.DIODE(\core_0.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__D (.DIODE(\core_0.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__A1 (.DIODE(\core_0.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__B2 (.DIODE(\core_0.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__D (.DIODE(\core_0.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A (.DIODE(\core_0.execute.rf.reg_outputs[6][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__D (.DIODE(\core_0.execute.rf.reg_outputs[6][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__D (.DIODE(\core_0.execute.rf.reg_outputs[6][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A (.DIODE(\core_0.execute.rf.reg_outputs[6][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__D (.DIODE(\core_0.execute.rf.reg_outputs[6][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A (.DIODE(\core_0.execute.rf.reg_outputs[6][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A (.DIODE(\core_0.execute.rf.reg_outputs[6][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__A (.DIODE(\core_0.execute.rf.reg_outputs[6][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__D (.DIODE(\core_0.execute.rf.reg_outputs[6][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A1 (.DIODE(\core_0.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__B2 (.DIODE(\core_0.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__B2 (.DIODE(\core_0.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__A (.DIODE(\core_0.execute.rf.reg_outputs[7][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A (.DIODE(\core_0.execute.rf.reg_outputs[7][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A (.DIODE(\core_0.execute.rf.reg_outputs[7][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A1 (.DIODE(\core_0.execute.rf.reg_outputs[7][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__B2 (.DIODE(\core_0.execute.rf.reg_outputs[7][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A (.DIODE(\core_0.execute.rf.reg_outputs[7][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A1 (.DIODE(\core_0.execute.rf.reg_outputs[7][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__B2 (.DIODE(\core_0.execute.rf.reg_outputs[7][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__A (.DIODE(\core_0.execute.rf.reg_outputs[7][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A1 (.DIODE(\core_0.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A1 (.DIODE(\core_0.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A (.DIODE(\core_0.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A1 (.DIODE(\core_0.execute.rf.reg_outputs[7][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A1 (.DIODE(\core_0.execute.rf.reg_outputs[7][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A1 (.DIODE(\core_0.execute.rf.reg_outputs[7][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A (.DIODE(\core_0.execute.rf.reg_outputs[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A (.DIODE(\core_0.execute.rf.reg_outputs[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A (.DIODE(\core_0.execute.rf.reg_outputs[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A (.DIODE(\core_0.execute.rf.reg_outputs[7][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A (.DIODE(\core_0.execute.rf.reg_outputs[7][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A1 (.DIODE(\core_0.execute.rf.reg_outputs[7][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A (.DIODE(\core_0.execute.rf.reg_outputs[7][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__A (.DIODE(\core_0.execute.rf.reg_outputs[7][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A (.DIODE(\core_0.execute.rf.reg_outputs[7][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A1 (.DIODE(\core_0.execute.rf.reg_outputs[7][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__A1 (.DIODE(\core_0.execute.rf.reg_outputs[7][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A (.DIODE(\core_0.execute.rf.reg_outputs[7][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A1 (.DIODE(\core_0.execute.rf.reg_outputs[7][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__B2 (.DIODE(\core_0.execute.rf.reg_outputs[7][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A (.DIODE(\core_0.execute.rf.reg_outputs[7][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__B2 (.DIODE(\core_0.execute.sreg_irq_flags.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A1 (.DIODE(\core_0.execute.sreg_irq_flags.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A (.DIODE(\core_0.execute.sreg_irq_flags.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A1 (.DIODE(\core_0.execute.sreg_irq_flags.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__B2 (.DIODE(\core_0.execute.sreg_irq_flags.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A1 (.DIODE(\core_0.execute.sreg_irq_flags.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A (.DIODE(\core_0.execute.sreg_irq_pc.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A (.DIODE(\core_0.execute.sreg_irq_pc.o_d[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A (.DIODE(\core_0.execute.sreg_irq_pc.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A (.DIODE(\core_0.execute.sreg_irq_pc.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A (.DIODE(\core_0.execute.sreg_irq_pc.o_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A (.DIODE(\core_0.execute.sreg_irq_pc.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A0 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A (.DIODE(\core_0.execute.sreg_irq_pc.o_d[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A1 (.DIODE(\core_0.execute.sreg_irq_pc.o_d[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A1 (.DIODE(\core_0.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__B2 (.DIODE(\core_0.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A (.DIODE(\core_0.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A1 (.DIODE(\core_0.execute.sreg_scratch.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__B2 (.DIODE(\core_0.execute.sreg_scratch.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A1 (.DIODE(\core_0.execute.sreg_scratch.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__B2 (.DIODE(\core_0.execute.sreg_scratch.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__A1 (.DIODE(\core_0.execute.sreg_scratch.o_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__B2 (.DIODE(\core_0.execute.sreg_scratch.o_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A1 (.DIODE(\core_0.execute.sreg_scratch.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__B2 (.DIODE(\core_0.execute.sreg_scratch.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A1 (.DIODE(\core_0.execute.sreg_scratch.o_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B2 (.DIODE(\core_0.execute.sreg_scratch.o_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_i_clk_A (.DIODE(i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(i_core_int_sreg[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(i_core_int_sreg[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(i_core_int_sreg[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(i_core_int_sreg[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(i_core_int_sreg[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(i_core_int_sreg[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(i_core_int_sreg[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(i_core_int_sreg[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(i_core_int_sreg[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(i_core_int_sreg[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(i_core_int_sreg[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(i_core_int_sreg[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(i_core_int_sreg[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(i_core_int_sreg[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(i_core_int_sreg[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(i_core_int_sreg[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(i_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(i_irq));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(i_mc_core_int));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(i_mem_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(i_mem_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(i_mem_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(i_mem_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(i_mem_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(i_mem_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(i_mem_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(i_mem_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(i_mem_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(i_mem_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(i_mem_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(i_mem_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(i_mem_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(i_mem_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(i_mem_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(i_mem_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(i_mem_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(i_mem_exception));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(i_req_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(i_req_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(i_req_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(i_req_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(i_req_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(i_req_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(i_req_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(i_req_data[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(i_req_data[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(i_req_data[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(i_req_data[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(i_req_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(i_req_data[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(i_req_data[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(i_req_data[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(i_req_data[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(i_req_data[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(i_req_data[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(i_req_data[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(i_req_data[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(i_req_data[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(i_req_data[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(i_req_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(i_req_data[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(i_req_data[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(i_req_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(i_req_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(i_req_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(i_req_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(i_req_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(i_req_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(i_req_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(i_req_data_valid));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(i_rst));
 sky130_fd_sc_hd__diode_2 ANTENNA__7289__CLK (.DIODE(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7291__CLK (.DIODE(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__CLK (.DIODE(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7293__CLK (.DIODE(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7296__CLK (.DIODE(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7295__CLK (.DIODE(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__B2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__B2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__B2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__B2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__B2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__B2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__A1_N (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A1_N (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A1_N (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A1_N (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__A0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A0 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A0 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__A0 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A0 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A0 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A0 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__D_N (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__C (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A1_N (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__A1_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__A1_N (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__A1_N (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A1_N (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__A1_N (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__A1_N (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__B2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A_N (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__S (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_output173_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_output176_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_output178_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A_N (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A0 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A_N (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_output179_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__C (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_output180_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_output181_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_output182_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__A0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__D (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_output183_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__C (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_output184_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_output185_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__C (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A_N (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_output186_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A_N (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A_N (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__A0 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_output187_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__D (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__D (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A_N (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A0 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__A0 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_output188_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__A0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_output189_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__A0 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_output190_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__D (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_output191_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__A0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__C (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_output192_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A_N (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A_N (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__B_N (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__B2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_output195_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_output196_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_output197_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_output198_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_output199_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__B1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_output200_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_output201_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_output202_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_output203_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_output204_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_output205_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_output206_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__A0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_output207_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_output208_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_output209_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_output210_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7258__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7251__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7254__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7256__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7240__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7242__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7236__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7241__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7235__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7191__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7189__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7190__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7199__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7200__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7174__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7232__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7203__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7204__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7171__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7183__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7186__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7201__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7170__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7233__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7217__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7234__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7218__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7215__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7231__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7263__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7250__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7248__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7147__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7244__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7246__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7243__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7265__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7262__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7268__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7146__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7196__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7279__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7198__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7212__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7213__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7230__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7166__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7270__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7269__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7266__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7282__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7261__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7260__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7259__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7281__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7278__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7020__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7019__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7022__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6978__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7016__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7018__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6988__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7139__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7120__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7301__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7153__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7371__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7360__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7369__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7370__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7372__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7368__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6881__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7348__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7350__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7349__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7347__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7353__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7352__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7374__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7373__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7364__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7365__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7133__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7327__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7329__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7330__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7351__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7321__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7322__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7320__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7319__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7324__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7323__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7325__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7326__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7318__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7332__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7331__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7343__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7345__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7344__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7342__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7380__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7376__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7341__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7340__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7355__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7356__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7359__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7358__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7377__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7354__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7339__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7338__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7378__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7098__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7357__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7388__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7381__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7382__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7093__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7362__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7396__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7333__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7392__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7395__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7366__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7361__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7375__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7363__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7367__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7335__CLK (.DIODE(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__CLK (.DIODE(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__CLK (.DIODE(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7336__CLK (.DIODE(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7334__CLK (.DIODE(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__CLK (.DIODE(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__CLK (.DIODE(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__CLK (.DIODE(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__CLK (.DIODE(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__CLK (.DIODE(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7316__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7061__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7384__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7383__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7385__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7300__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7306__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7309__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7310__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7294__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7297__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7299__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7298__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7054__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7305__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_i_clk_A (.DIODE(clknet_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_i_clk_A (.DIODE(clknet_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_i_clk_A (.DIODE(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_i_clk_A (.DIODE(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_i_clk_A (.DIODE(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_i_clk_A (.DIODE(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_1_0_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_286_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_286_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_286_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_286_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_288_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_290_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_290_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_841 ();
 assign o_mem_addr_high[7] = net211;
endmodule

