// This is the unpowered netlist.
module interconnect_outer (inner_clock,
    inner_disable,
    inner_embed_mode,
    inner_ext_irq,
    inner_reset,
    inner_wb_4_burst,
    inner_wb_8_burst,
    inner_wb_ack,
    inner_wb_cyc,
    inner_wb_err,
    inner_wb_stb,
    inner_wb_we,
    iram1_clk,
    iram1_csb,
    iram_clk,
    iram_csb,
    iram_we,
    mgt_wb_ack_o,
    mgt_wb_clk_i,
    mgt_wb_cyc_i,
    mgt_wb_rst_i,
    mgt_wb_stb_i,
    mgt_wb_we_i,
    user_clock2,
    inner_wb_adr,
    inner_wb_i_dat,
    inner_wb_o_dat,
    inner_wb_sel,
    iram1_addr,
    iram1_dout,
    iram_addr,
    iram_i_data,
    iram_o_data,
    iram_w_mask,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    m_io_in,
    m_io_oeb,
    m_io_out,
    mgt_wb_adr_i,
    mgt_wb_dat_i,
    mgt_wb_dat_o,
    mgt_wb_sel_i);
 output inner_clock;
 output inner_disable;
 output inner_embed_mode;
 output inner_ext_irq;
 output inner_reset;
 input inner_wb_4_burst;
 input inner_wb_8_burst;
 output inner_wb_ack;
 input inner_wb_cyc;
 output inner_wb_err;
 input inner_wb_stb;
 input inner_wb_we;
 input iram1_clk;
 input iram1_csb;
 output iram_clk;
 output iram_csb;
 output iram_we;
 output mgt_wb_ack_o;
 input mgt_wb_clk_i;
 input mgt_wb_cyc_i;
 input mgt_wb_rst_i;
 input mgt_wb_stb_i;
 input mgt_wb_we_i;
 input user_clock2;
 input [23:0] inner_wb_adr;
 output [15:0] inner_wb_i_dat;
 input [15:0] inner_wb_o_dat;
 input [1:0] inner_wb_sel;
 output [7:0] iram1_addr;
 input [31:0] iram1_dout;
 output [7:0] iram_addr;
 output [31:0] iram_i_data;
 input [31:0] iram_o_data;
 output [3:0] iram_w_mask;
 output [2:0] irq;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [37:0] m_io_in;
 output [37:0] m_io_oeb;
 output [37:0] m_io_out;
 input [31:0] mgt_wb_adr_i;
 input [31:0] mgt_wb_dat_i;
 output [31:0] mgt_wb_dat_o;
 input [3:0] mgt_wb_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire net206;
 wire net207;
 wire \clk_div.clock_sel ;
 wire \clk_div.clock_sel_r ;
 wire \clk_div.cnt[0] ;
 wire \clk_div.cnt[10] ;
 wire \clk_div.cnt[11] ;
 wire \clk_div.cnt[12] ;
 wire \clk_div.cnt[13] ;
 wire \clk_div.cnt[14] ;
 wire \clk_div.cnt[15] ;
 wire \clk_div.cnt[1] ;
 wire \clk_div.cnt[2] ;
 wire \clk_div.cnt[3] ;
 wire \clk_div.cnt[4] ;
 wire \clk_div.cnt[5] ;
 wire \clk_div.cnt[6] ;
 wire \clk_div.cnt[7] ;
 wire \clk_div.cnt[8] ;
 wire \clk_div.cnt[9] ;
 wire \clk_div.curr_div[0] ;
 wire \clk_div.curr_div[1] ;
 wire \clk_div.curr_div[2] ;
 wire \clk_div.curr_div[3] ;
 wire \clk_div.next_div_buff[0] ;
 wire \clk_div.next_div_buff[1] ;
 wire \clk_div.next_div_buff[2] ;
 wire \clk_div.next_div_buff[3] ;
 wire \clk_div.next_div_val ;
 wire \clk_div.res_clk ;
 wire \disable_s_ff[0] ;
 wire \embed_s_ff[0] ;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net414;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire iram_wb_ack;
 wire net236;
 wire net237;
 wire net238;
 wire \irq_s_ff[0] ;
 wire net239;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net249;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net250;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net240;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net241;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net242;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net243;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net244;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net245;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net246;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net247;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net248;
 wire \m_arbiter.i_wb0_cyc ;
 wire \m_arbiter.o_sel_sig ;
 wire \m_arbiter.wb0_adr[0] ;
 wire \m_arbiter.wb0_adr[10] ;
 wire \m_arbiter.wb0_adr[11] ;
 wire \m_arbiter.wb0_adr[12] ;
 wire \m_arbiter.wb0_adr[13] ;
 wire \m_arbiter.wb0_adr[14] ;
 wire \m_arbiter.wb0_adr[15] ;
 wire \m_arbiter.wb0_adr[16] ;
 wire \m_arbiter.wb0_adr[17] ;
 wire \m_arbiter.wb0_adr[18] ;
 wire \m_arbiter.wb0_adr[19] ;
 wire \m_arbiter.wb0_adr[1] ;
 wire \m_arbiter.wb0_adr[20] ;
 wire \m_arbiter.wb0_adr[21] ;
 wire \m_arbiter.wb0_adr[22] ;
 wire \m_arbiter.wb0_adr[23] ;
 wire \m_arbiter.wb0_adr[2] ;
 wire \m_arbiter.wb0_adr[3] ;
 wire \m_arbiter.wb0_adr[4] ;
 wire \m_arbiter.wb0_adr[5] ;
 wire \m_arbiter.wb0_adr[6] ;
 wire \m_arbiter.wb0_adr[7] ;
 wire \m_arbiter.wb0_adr[8] ;
 wire \m_arbiter.wb0_adr[9] ;
 wire \m_arbiter.wb0_o_dat[0] ;
 wire \m_arbiter.wb0_o_dat[10] ;
 wire \m_arbiter.wb0_o_dat[11] ;
 wire \m_arbiter.wb0_o_dat[12] ;
 wire \m_arbiter.wb0_o_dat[13] ;
 wire \m_arbiter.wb0_o_dat[14] ;
 wire \m_arbiter.wb0_o_dat[15] ;
 wire \m_arbiter.wb0_o_dat[1] ;
 wire \m_arbiter.wb0_o_dat[2] ;
 wire \m_arbiter.wb0_o_dat[3] ;
 wire \m_arbiter.wb0_o_dat[4] ;
 wire \m_arbiter.wb0_o_dat[5] ;
 wire \m_arbiter.wb0_o_dat[6] ;
 wire \m_arbiter.wb0_o_dat[7] ;
 wire \m_arbiter.wb0_o_dat[8] ;
 wire \m_arbiter.wb0_o_dat[9] ;
 wire \m_arbiter.wb0_we ;
 wire net415;
 wire net416;
 wire net369;
 wire net370;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net371;
 wire net372;
 wire net367;
 wire net368;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire clknet_leaf_0_user_clock2;
 wire net381;
 wire net382;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net383;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net384;
 wire net412;
 wire net413;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire \rst_cw_sync.reset_sync_ff[0] ;
 wire \rst_soc_sync.reset_sync_ff[0] ;
 wire \split_s_ff[0] ;
 wire \sspi.bit_cnt[0] ;
 wire \sspi.bit_cnt[1] ;
 wire \sspi.bit_cnt[2] ;
 wire \sspi.bit_cnt[3] ;
 wire \sspi.bit_cnt[4] ;
 wire \sspi.req_addr[0] ;
 wire \sspi.req_addr[10] ;
 wire \sspi.req_addr[11] ;
 wire \sspi.req_addr[12] ;
 wire \sspi.req_addr[13] ;
 wire \sspi.req_addr[14] ;
 wire \sspi.req_addr[15] ;
 wire \sspi.req_addr[16] ;
 wire \sspi.req_addr[17] ;
 wire \sspi.req_addr[18] ;
 wire \sspi.req_addr[19] ;
 wire \sspi.req_addr[1] ;
 wire \sspi.req_addr[20] ;
 wire \sspi.req_addr[21] ;
 wire \sspi.req_addr[22] ;
 wire \sspi.req_addr[23] ;
 wire \sspi.req_addr[2] ;
 wire \sspi.req_addr[3] ;
 wire \sspi.req_addr[4] ;
 wire \sspi.req_addr[5] ;
 wire \sspi.req_addr[6] ;
 wire \sspi.req_addr[7] ;
 wire \sspi.req_addr[8] ;
 wire \sspi.req_addr[9] ;
 wire \sspi.req_data[0] ;
 wire \sspi.req_data[10] ;
 wire \sspi.req_data[11] ;
 wire \sspi.req_data[12] ;
 wire \sspi.req_data[13] ;
 wire \sspi.req_data[14] ;
 wire \sspi.req_data[15] ;
 wire \sspi.req_data[1] ;
 wire \sspi.req_data[2] ;
 wire \sspi.req_data[3] ;
 wire \sspi.req_data[4] ;
 wire \sspi.req_data[5] ;
 wire \sspi.req_data[6] ;
 wire \sspi.req_data[7] ;
 wire \sspi.req_data[8] ;
 wire \sspi.req_data[9] ;
 wire \sspi.res_data[0] ;
 wire \sspi.res_data[10] ;
 wire \sspi.res_data[11] ;
 wire \sspi.res_data[12] ;
 wire \sspi.res_data[13] ;
 wire \sspi.res_data[14] ;
 wire \sspi.res_data[15] ;
 wire \sspi.res_data[1] ;
 wire \sspi.res_data[2] ;
 wire \sspi.res_data[3] ;
 wire \sspi.res_data[4] ;
 wire \sspi.res_data[5] ;
 wire \sspi.res_data[6] ;
 wire \sspi.res_data[7] ;
 wire \sspi.res_data[8] ;
 wire \sspi.res_data[9] ;
 wire \sspi.resp_err ;
 wire \sspi.state[0] ;
 wire \sspi.state[1] ;
 wire \sspi.state[2] ;
 wire \sspi.state[3] ;
 wire \sspi.state[4] ;
 wire \sspi.state[5] ;
 wire \sspi.state[6] ;
 wire \sspi.state[7] ;
 wire \sspi.sy_clk[0] ;
 wire \sspi.sy_clk[1] ;
 wire \sspi.sy_clk[2] ;
 wire \wb_compressor.burst_cnt[0] ;
 wire \wb_compressor.burst_cnt[1] ;
 wire \wb_compressor.burst_cnt[2] ;
 wire \wb_compressor.burst_end[0] ;
 wire \wb_compressor.burst_end[2] ;
 wire \wb_compressor.l_we ;
 wire \wb_compressor.state[0] ;
 wire \wb_compressor.state[1] ;
 wire \wb_compressor.state[2] ;
 wire \wb_compressor.state[3] ;
 wire \wb_compressor.state[4] ;
 wire \wb_compressor.state[5] ;
 wire \wb_compressor.state[6] ;
 wire \wb_compressor.wb_ack ;
 wire \wb_compressor.wb_err ;
 wire \wb_compressor.wb_i_dat[0] ;
 wire \wb_compressor.wb_i_dat[10] ;
 wire \wb_compressor.wb_i_dat[11] ;
 wire \wb_compressor.wb_i_dat[12] ;
 wire \wb_compressor.wb_i_dat[13] ;
 wire \wb_compressor.wb_i_dat[14] ;
 wire \wb_compressor.wb_i_dat[15] ;
 wire \wb_compressor.wb_i_dat[1] ;
 wire \wb_compressor.wb_i_dat[2] ;
 wire \wb_compressor.wb_i_dat[3] ;
 wire \wb_compressor.wb_i_dat[4] ;
 wire \wb_compressor.wb_i_dat[5] ;
 wire \wb_compressor.wb_i_dat[6] ;
 wire \wb_compressor.wb_i_dat[7] ;
 wire \wb_compressor.wb_i_dat[8] ;
 wire \wb_compressor.wb_i_dat[9] ;
 wire \wb_cross_clk.ack_next_hold ;
 wire \wb_cross_clk.ack_xor_flag ;
 wire \wb_cross_clk.err_xor_flag ;
 wire \wb_cross_clk.m_burst_cnt[0] ;
 wire \wb_cross_clk.m_burst_cnt[1] ;
 wire \wb_cross_clk.m_burst_cnt[2] ;
 wire \wb_cross_clk.m_burst_cnt[3] ;
 wire \wb_cross_clk.m_new_req_flag ;
 wire \wb_cross_clk.m_s_sync.d_data[0] ;
 wire \wb_cross_clk.m_s_sync.d_data[10] ;
 wire \wb_cross_clk.m_s_sync.d_data[11] ;
 wire \wb_cross_clk.m_s_sync.d_data[12] ;
 wire \wb_cross_clk.m_s_sync.d_data[13] ;
 wire \wb_cross_clk.m_s_sync.d_data[14] ;
 wire \wb_cross_clk.m_s_sync.d_data[15] ;
 wire \wb_cross_clk.m_s_sync.d_data[16] ;
 wire \wb_cross_clk.m_s_sync.d_data[17] ;
 wire \wb_cross_clk.m_s_sync.d_data[18] ;
 wire \wb_cross_clk.m_s_sync.d_data[19] ;
 wire \wb_cross_clk.m_s_sync.d_data[1] ;
 wire \wb_cross_clk.m_s_sync.d_data[20] ;
 wire \wb_cross_clk.m_s_sync.d_data[21] ;
 wire \wb_cross_clk.m_s_sync.d_data[22] ;
 wire \wb_cross_clk.m_s_sync.d_data[23] ;
 wire \wb_cross_clk.m_s_sync.d_data[24] ;
 wire \wb_cross_clk.m_s_sync.d_data[25] ;
 wire \wb_cross_clk.m_s_sync.d_data[26] ;
 wire \wb_cross_clk.m_s_sync.d_data[27] ;
 wire \wb_cross_clk.m_s_sync.d_data[28] ;
 wire \wb_cross_clk.m_s_sync.d_data[29] ;
 wire \wb_cross_clk.m_s_sync.d_data[2] ;
 wire \wb_cross_clk.m_s_sync.d_data[30] ;
 wire \wb_cross_clk.m_s_sync.d_data[31] ;
 wire \wb_cross_clk.m_s_sync.d_data[32] ;
 wire \wb_cross_clk.m_s_sync.d_data[33] ;
 wire \wb_cross_clk.m_s_sync.d_data[34] ;
 wire \wb_cross_clk.m_s_sync.d_data[35] ;
 wire \wb_cross_clk.m_s_sync.d_data[36] ;
 wire \wb_cross_clk.m_s_sync.d_data[37] ;
 wire \wb_cross_clk.m_s_sync.d_data[38] ;
 wire \wb_cross_clk.m_s_sync.d_data[39] ;
 wire \wb_cross_clk.m_s_sync.d_data[3] ;
 wire \wb_cross_clk.m_s_sync.d_data[40] ;
 wire \wb_cross_clk.m_s_sync.d_data[41] ;
 wire \wb_cross_clk.m_s_sync.d_data[42] ;
 wire \wb_cross_clk.m_s_sync.d_data[43] ;
 wire \wb_cross_clk.m_s_sync.d_data[44] ;
 wire \wb_cross_clk.m_s_sync.d_data[45] ;
 wire \wb_cross_clk.m_s_sync.d_data[46] ;
 wire \wb_cross_clk.m_s_sync.d_data[4] ;
 wire \wb_cross_clk.m_s_sync.d_data[5] ;
 wire \wb_cross_clk.m_s_sync.d_data[6] ;
 wire \wb_cross_clk.m_s_sync.d_data[7] ;
 wire \wb_cross_clk.m_s_sync.d_data[8] ;
 wire \wb_cross_clk.m_s_sync.d_data[9] ;
 wire \wb_cross_clk.m_s_sync.d_xfer_xor_sync[0] ;
 wire \wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ;
 wire \wb_cross_clk.m_s_sync.d_xfer_xor_sync[2] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[0] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[10] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[11] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[12] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[13] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[14] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[15] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[16] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[17] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[18] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[19] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[1] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[20] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[21] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[22] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[23] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[24] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[25] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[26] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[27] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[28] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[29] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[2] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[30] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[31] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[32] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[33] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[34] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[35] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[36] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[37] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[38] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[39] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[3] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[40] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[41] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[42] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[43] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[44] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[45] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[46] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[4] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[5] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[6] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[7] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[8] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[9] ;
 wire \wb_cross_clk.m_s_sync.s_xfer_xor_flag ;
 wire \wb_cross_clk.m_wb_i_dat[0] ;
 wire \wb_cross_clk.m_wb_i_dat[10] ;
 wire \wb_cross_clk.m_wb_i_dat[11] ;
 wire \wb_cross_clk.m_wb_i_dat[12] ;
 wire \wb_cross_clk.m_wb_i_dat[13] ;
 wire \wb_cross_clk.m_wb_i_dat[14] ;
 wire \wb_cross_clk.m_wb_i_dat[15] ;
 wire \wb_cross_clk.m_wb_i_dat[1] ;
 wire \wb_cross_clk.m_wb_i_dat[2] ;
 wire \wb_cross_clk.m_wb_i_dat[3] ;
 wire \wb_cross_clk.m_wb_i_dat[4] ;
 wire \wb_cross_clk.m_wb_i_dat[5] ;
 wire \wb_cross_clk.m_wb_i_dat[6] ;
 wire \wb_cross_clk.m_wb_i_dat[7] ;
 wire \wb_cross_clk.m_wb_i_dat[8] ;
 wire \wb_cross_clk.m_wb_i_dat[9] ;
 wire \wb_cross_clk.msy_xor_ack ;
 wire \wb_cross_clk.msy_xor_err ;
 wire \wb_cross_clk.prev_ack ;
 wire \wb_cross_clk.prev_stb ;
 wire \wb_cross_clk.prev_xor_ack ;
 wire \wb_cross_clk.prev_xor_err ;
 wire \wb_cross_clk.prev_xor_newreq ;
 wire \wb_cross_clk.s_burst_cnt[0] ;
 wire \wb_cross_clk.s_burst_cnt[1] ;
 wire \wb_cross_clk.s_burst_cnt[2] ;
 wire \wb_cross_clk.s_burst_cnt[3] ;
 wire \wb_cross_clk.s_m_sync.d_xfer_xor_sync[0] ;
 wire \wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ;
 wire \wb_cross_clk.s_m_sync.d_xfer_xor_sync[2] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[0] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[10] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[11] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[12] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[13] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[14] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[15] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[16] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[17] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[1] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[2] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[3] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[4] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[5] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[6] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[7] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[8] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[9] ;
 wire \wb_cross_clk.s_m_sync.s_xfer_xor_flag ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire clknet_leaf_1_user_clock2;
 wire clknet_leaf_2_user_clock2;
 wire clknet_leaf_3_user_clock2;
 wire clknet_leaf_4_user_clock2;
 wire clknet_leaf_5_user_clock2;
 wire clknet_leaf_6_user_clock2;
 wire clknet_leaf_7_user_clock2;
 wire clknet_leaf_8_user_clock2;
 wire clknet_leaf_9_user_clock2;
 wire clknet_leaf_10_user_clock2;
 wire clknet_leaf_11_user_clock2;
 wire clknet_leaf_12_user_clock2;
 wire clknet_leaf_13_user_clock2;
 wire clknet_leaf_14_user_clock2;
 wire clknet_leaf_15_user_clock2;
 wire clknet_leaf_16_user_clock2;
 wire clknet_leaf_17_user_clock2;
 wire clknet_leaf_18_user_clock2;
 wire clknet_leaf_19_user_clock2;
 wire clknet_leaf_20_user_clock2;
 wire clknet_leaf_22_user_clock2;
 wire clknet_leaf_23_user_clock2;
 wire clknet_leaf_24_user_clock2;
 wire clknet_leaf_25_user_clock2;
 wire clknet_leaf_26_user_clock2;
 wire clknet_leaf_27_user_clock2;
 wire clknet_leaf_28_user_clock2;
 wire clknet_leaf_29_user_clock2;
 wire clknet_leaf_30_user_clock2;
 wire clknet_leaf_31_user_clock2;
 wire clknet_leaf_32_user_clock2;
 wire clknet_leaf_33_user_clock2;
 wire clknet_leaf_34_user_clock2;
 wire clknet_leaf_36_user_clock2;
 wire clknet_0_user_clock2;
 wire clknet_2_0__leaf_user_clock2;
 wire clknet_2_1__leaf_user_clock2;
 wire clknet_2_2__leaf_user_clock2;
 wire clknet_2_3__leaf_user_clock2;
 wire clknet_opt_1_0_user_clock2;
 wire clknet_opt_2_0_user_clock2;
 wire clknet_0_net190;
 wire clknet_4_0_0_net190;
 wire clknet_4_1_0_net190;
 wire clknet_4_2_0_net190;
 wire clknet_4_3_0_net190;
 wire clknet_4_4_0_net190;
 wire clknet_4_5_0_net190;
 wire clknet_4_6_0_net190;
 wire clknet_4_7_0_net190;
 wire clknet_4_8_0_net190;
 wire clknet_4_9_0_net190;
 wire clknet_4_10_0_net190;
 wire clknet_4_11_0_net190;
 wire clknet_4_12_0_net190;
 wire clknet_4_13_0_net190;
 wire clknet_4_14_0_net190;
 wire clknet_4_15_0_net190;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;

 sky130_fd_sc_hd__buf_4 _1329_ (.A(\m_arbiter.o_sel_sig ),
    .X(_1224_));
 sky130_fd_sc_hd__buf_4 _1330_ (.A(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__mux2_1 _1331_ (.A0(net640),
    .A1(net41),
    .S(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_4 _1332_ (.A(_1226_),
    .X(net144));
 sky130_fd_sc_hd__mux2_1 _1333_ (.A0(net647),
    .A1(net40),
    .S(_1225_),
    .X(_1227_));
 sky130_fd_sc_hd__buf_4 _1334_ (.A(net648),
    .X(net143));
 sky130_fd_sc_hd__mux2_1 _1335_ (.A0(net678),
    .A1(net39),
    .S(_1224_),
    .X(_1228_));
 sky130_fd_sc_hd__buf_4 _1336_ (.A(net679),
    .X(net142));
 sky130_fd_sc_hd__buf_4 _1337_ (.A(_1224_),
    .X(_1229_));
 sky130_fd_sc_hd__mux2_1 _1338_ (.A0(net652),
    .A1(net38),
    .S(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__buf_4 _1339_ (.A(_1230_),
    .X(net141));
 sky130_fd_sc_hd__mux2_1 _1340_ (.A0(net594),
    .A1(net37),
    .S(_1229_),
    .X(_1231_));
 sky130_fd_sc_hd__buf_4 _1341_ (.A(net595),
    .X(net140));
 sky130_fd_sc_hd__mux2_1 _1342_ (.A0(net615),
    .A1(net36),
    .S(_1225_),
    .X(_1232_));
 sky130_fd_sc_hd__buf_4 _1343_ (.A(net616),
    .X(net139));
 sky130_fd_sc_hd__mux2_1 _1344_ (.A0(\m_arbiter.wb0_o_dat[1] ),
    .A1(net35),
    .S(_1229_),
    .X(_1233_));
 sky130_fd_sc_hd__buf_4 _1345_ (.A(_1233_),
    .X(net138));
 sky130_fd_sc_hd__mux2_1 _1346_ (.A0(\m_arbiter.wb0_o_dat[0] ),
    .A1(net28),
    .S(_1224_),
    .X(_1234_));
 sky130_fd_sc_hd__buf_4 _1347_ (.A(_1234_),
    .X(net131));
 sky130_fd_sc_hd__buf_4 _1348_ (.A(\m_arbiter.o_sel_sig ),
    .X(_1235_));
 sky130_fd_sc_hd__mux2_1 _1349_ (.A0(\m_arbiter.wb0_adr[3] ),
    .A1(net20),
    .S(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__clkbuf_4 _1350_ (.A(_1236_),
    .X(net125));
 sky130_fd_sc_hd__mux2_1 _1351_ (.A0(\m_arbiter.wb0_adr[2] ),
    .A1(net19),
    .S(_1235_),
    .X(_1237_));
 sky130_fd_sc_hd__clkbuf_4 _1352_ (.A(_1237_),
    .X(net124));
 sky130_fd_sc_hd__mux2_1 _1353_ (.A0(net625),
    .A1(net14),
    .S(_1235_),
    .X(_1238_));
 sky130_fd_sc_hd__buf_4 _1354_ (.A(net626),
    .X(net123));
 sky130_fd_sc_hd__buf_4 _1355_ (.A(\m_arbiter.o_sel_sig ),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_1 _1356_ (.A0(net657),
    .A1(net3),
    .S(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__clkbuf_4 _1357_ (.A(net658),
    .X(net122));
 sky130_fd_sc_hd__mux2_1 _1358_ (.A0(\m_arbiter.wb0_adr[7] ),
    .A1(net24),
    .S(\m_arbiter.o_sel_sig ),
    .X(_1241_));
 sky130_fd_sc_hd__clkbuf_2 _1359_ (.A(_1241_),
    .X(net129));
 sky130_fd_sc_hd__mux2_1 _1360_ (.A0(\m_arbiter.wb0_adr[6] ),
    .A1(net23),
    .S(_1235_),
    .X(_1242_));
 sky130_fd_sc_hd__buf_2 _1361_ (.A(_1242_),
    .X(net128));
 sky130_fd_sc_hd__mux2_1 _1362_ (.A0(\m_arbiter.wb0_adr[5] ),
    .A1(net22),
    .S(_1235_),
    .X(_1243_));
 sky130_fd_sc_hd__buf_2 _1363_ (.A(_1243_),
    .X(net127));
 sky130_fd_sc_hd__mux2_1 _1364_ (.A0(\m_arbiter.wb0_adr[4] ),
    .A1(net21),
    .S(_1224_),
    .X(_1244_));
 sky130_fd_sc_hd__clkbuf_4 _1365_ (.A(_1244_),
    .X(net126));
 sky130_fd_sc_hd__or2_1 _1366_ (.A(net125),
    .B(net124),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_1 _1367_ (.A0(net582),
    .A1(net12),
    .S(_1235_),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_2 _1368_ (.A0(net620),
    .A1(net11),
    .S(_1235_),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _1369_ (.A0(net587),
    .A1(net13),
    .S(_1239_),
    .X(_1248_));
 sky130_fd_sc_hd__mux2_1 _1370_ (.A0(net605),
    .A1(net10),
    .S(_1239_),
    .X(_1249_));
 sky130_fd_sc_hd__or4_2 _1371_ (.A(_1246_),
    .B(_1247_),
    .C(_1248_),
    .D(_1249_),
    .X(_1250_));
 sky130_fd_sc_hd__mux2_2 _1372_ (.A0(\m_arbiter.wb0_adr[23] ),
    .A1(net18),
    .S(_1235_),
    .X(_1251_));
 sky130_fd_sc_hd__mux2_2 _1373_ (.A0(net610),
    .A1(net15),
    .S(_1235_),
    .X(_1252_));
 sky130_fd_sc_hd__mux2_4 _1374_ (.A0(net634),
    .A1(net16),
    .S(_1235_),
    .X(_1253_));
 sky130_fd_sc_hd__mux2_2 _1375_ (.A0(net630),
    .A1(net17),
    .S(_1239_),
    .X(_1254_));
 sky130_fd_sc_hd__or4_1 _1376_ (.A(_1251_),
    .B(_1252_),
    .C(_1253_),
    .D(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__or3_2 _1377_ (.A(_1245_),
    .B(_1250_),
    .C(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__mux2_2 _1378_ (.A0(\m_arbiter.wb0_adr[12] ),
    .A1(net6),
    .S(_1224_),
    .X(_1257_));
 sky130_fd_sc_hd__inv_2 _1379_ (.A(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__mux2_2 _1380_ (.A0(net836),
    .A1(net7),
    .S(_1239_),
    .X(_1259_));
 sky130_fd_sc_hd__mux2_2 _1381_ (.A0(net600),
    .A1(net8),
    .S(_1239_),
    .X(_1260_));
 sky130_fd_sc_hd__mux2_1 _1382_ (.A0(net577),
    .A1(net9),
    .S(_1224_),
    .X(_1261_));
 sky130_fd_sc_hd__or3_1 _1383_ (.A(_1259_),
    .B(_1260_),
    .C(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__mux2_2 _1384_ (.A0(\m_arbiter.wb0_adr[8] ),
    .A1(net25),
    .S(_1239_),
    .X(_1263_));
 sky130_fd_sc_hd__mux2_1 _1385_ (.A0(net818),
    .A1(net4),
    .S(_1239_),
    .X(_1264_));
 sky130_fd_sc_hd__mux2_2 _1386_ (.A0(\m_arbiter.wb0_adr[9] ),
    .A1(net26),
    .S(_1239_),
    .X(_1265_));
 sky130_fd_sc_hd__mux2_2 _1387_ (.A0(net741),
    .A1(net5),
    .S(_1239_),
    .X(_1266_));
 sky130_fd_sc_hd__or4_1 _1388_ (.A(_1263_),
    .B(_1264_),
    .C(_1265_),
    .D(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__or3_4 _1389_ (.A(_1258_),
    .B(_1262_),
    .C(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__or4b_1 _1390_ (.A(net129),
    .B(net128),
    .C(net127),
    .D_N(net126),
    .X(_1269_));
 sky130_fd_sc_hd__a2111o_1 _1391_ (.A1(net123),
    .A2(net122),
    .B1(_1256_),
    .C1(_1268_),
    .D1(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__and4_2 _1392_ (.A(_1246_),
    .B(_1247_),
    .C(_1248_),
    .D(_1254_),
    .X(_1271_));
 sky130_fd_sc_hd__and3_1 _1393_ (.A(_1257_),
    .B(_1265_),
    .C(_1266_),
    .X(_1272_));
 sky130_fd_sc_hd__and4b_1 _1394_ (.A_N(_1263_),
    .B(_1264_),
    .C(_1259_),
    .D(_1261_),
    .X(_1273_));
 sky130_fd_sc_hd__and4b_1 _1395_ (.A_N(_1251_),
    .B(_1252_),
    .C(_1249_),
    .D(_1260_),
    .X(_1274_));
 sky130_fd_sc_hd__and3_2 _1396_ (.A(_1272_),
    .B(_1273_),
    .C(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__a31oi_4 _1397_ (.A1(net635),
    .A2(_1271_),
    .A3(_1275_),
    .B1(net90),
    .Y(_1276_));
 sky130_fd_sc_hd__or3_1 _1398_ (.A(net129),
    .B(net128),
    .C(net127),
    .X(_1277_));
 sky130_fd_sc_hd__or2b_1 _1399_ (.A(net123),
    .B_N(net122),
    .X(_1278_));
 sky130_fd_sc_hd__or3_1 _1400_ (.A(net126),
    .B(_1277_),
    .C(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__or3_2 _1401_ (.A(_1256_),
    .B(_1268_),
    .C(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__or2b_1 _1402_ (.A(_1224_),
    .B_N(\m_arbiter.i_wb0_cyc ),
    .X(_1281_));
 sky130_fd_sc_hd__a21bo_1 _1403_ (.A1(_1224_),
    .A2(net46),
    .B1_N(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__nand2_1 _1404_ (.A(_1224_),
    .B(net27),
    .Y(_1283_));
 sky130_fd_sc_hd__a21oi_2 _1405_ (.A1(_1281_),
    .A2(_1283_),
    .B1(net103),
    .Y(_1284_));
 sky130_fd_sc_hd__and2_2 _1406_ (.A(_1282_),
    .B(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__and2b_1 _1407_ (.A_N(\wb_cross_clk.ack_next_hold ),
    .B(\wb_cross_clk.m_s_sync.d_data[46] ),
    .X(_1286_));
 sky130_fd_sc_hd__mux2_1 _1408_ (.A0(_1285_),
    .A1(_1286_),
    .S(net204),
    .X(_1287_));
 sky130_fd_sc_hd__and4_1 _1409_ (.A(_1270_),
    .B(net636),
    .C(_1280_),
    .D(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_4 _1410_ (.A(net637),
    .X(_1289_));
 sky130_fd_sc_hd__o21ai_4 _1411_ (.A1(net85),
    .A2(net84),
    .B1(_1289_),
    .Y(_1290_));
 sky130_fd_sc_hd__or2_1 _1412_ (.A(\wb_compressor.burst_end[2] ),
    .B(\wb_compressor.burst_cnt[2] ),
    .X(_1291_));
 sky130_fd_sc_hd__nand2_1 _1413_ (.A(\wb_compressor.burst_end[2] ),
    .B(\wb_compressor.burst_cnt[2] ),
    .Y(_1292_));
 sky130_fd_sc_hd__nand2_1 _1414_ (.A(\wb_compressor.burst_cnt[0] ),
    .B(\wb_compressor.burst_cnt[1] ),
    .Y(_1293_));
 sky130_fd_sc_hd__nor2_1 _1415_ (.A(\wb_compressor.burst_cnt[0] ),
    .B(\wb_compressor.burst_cnt[1] ),
    .Y(_1294_));
 sky130_fd_sc_hd__nor2_1 _1416_ (.A(\wb_compressor.burst_end[0] ),
    .B(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__a221o_1 _1417_ (.A1(_1291_),
    .A2(_1292_),
    .B1(_1293_),
    .B2(\wb_compressor.burst_end[0] ),
    .C1(_1295_),
    .X(_1296_));
 sky130_fd_sc_hd__o21ai_1 _1418_ (.A1(_1290_),
    .A2(_1296_),
    .B1(\wb_compressor.state[5] ),
    .Y(_1297_));
 sky130_fd_sc_hd__nand3b_1 _1419_ (.A_N(net575),
    .B(net84),
    .C(net690),
    .Y(_1298_));
 sky130_fd_sc_hd__a21oi_1 _1420_ (.A1(_1297_),
    .A2(_1298_),
    .B1(net201),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1421_ (.A(net201),
    .Y(_1299_));
 sky130_fd_sc_hd__buf_2 _1422_ (.A(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__inv_2 _1423_ (.A(_1290_),
    .Y(_1301_));
 sky130_fd_sc_hd__inv_2 _1424_ (.A(\wb_compressor.wb_ack ),
    .Y(_1302_));
 sky130_fd_sc_hd__a21boi_2 _1425_ (.A1(_1302_),
    .A2(_1289_),
    .B1_N(\wb_compressor.state[6] ),
    .Y(_1303_));
 sky130_fd_sc_hd__a31o_1 _1426_ (.A1(net957),
    .A2(_1301_),
    .A3(_1296_),
    .B1(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__and2_1 _1427_ (.A(_1300_),
    .B(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_1 _1428_ (.A(_1305_),
    .X(_0014_));
 sky130_fd_sc_hd__nand3_1 _1429_ (.A(_1302_),
    .B(net668),
    .C(_1289_),
    .Y(_1306_));
 sky130_fd_sc_hd__a32o_1 _1430_ (.A1(\wb_compressor.state[2] ),
    .A2(net84),
    .A3(net575),
    .B1(_1290_),
    .B2(\wb_compressor.state[4] ),
    .X(_1307_));
 sky130_fd_sc_hd__inv_2 _1431_ (.A(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__a21oi_1 _1432_ (.A1(net669),
    .A2(_1308_),
    .B1(net201),
    .Y(_0012_));
 sky130_fd_sc_hd__clkbuf_4 _1433_ (.A(\wb_compressor.state[3] ),
    .X(_1309_));
 sky130_fd_sc_hd__and2b_1 _1434_ (.A_N(net84),
    .B(net690),
    .X(_1310_));
 sky130_fd_sc_hd__clkbuf_4 _1435_ (.A(_1299_),
    .X(_1311_));
 sky130_fd_sc_hd__buf_2 _1436_ (.A(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__o21a_1 _1437_ (.A1(_1309_),
    .A2(_1310_),
    .B1(_1312_),
    .X(_0011_));
 sky130_fd_sc_hd__buf_4 _1438_ (.A(net204),
    .X(_1313_));
 sky130_fd_sc_hd__mux2_1 _1439_ (.A0(net621),
    .A1(\wb_cross_clk.m_s_sync.d_data[39] ),
    .S(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__mux2_1 _1440_ (.A0(_1251_),
    .A1(\wb_cross_clk.m_s_sync.d_data[45] ),
    .S(_1313_),
    .X(_1315_));
 sky130_fd_sc_hd__mux2_1 _1441_ (.A0(net635),
    .A1(\wb_cross_clk.m_s_sync.d_data[43] ),
    .S(_1313_),
    .X(_1316_));
 sky130_fd_sc_hd__or3_2 _1442_ (.A(_1314_),
    .B(_1315_),
    .C(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__mux2_1 _1443_ (.A0(net611),
    .A1(\wb_cross_clk.m_s_sync.d_data[42] ),
    .S(net204),
    .X(_1318_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(net578),
    .A1(\wb_cross_clk.m_s_sync.d_data[37] ),
    .S(net204),
    .X(_1319_));
 sky130_fd_sc_hd__mux2_1 _1445_ (.A0(net583),
    .A1(\wb_cross_clk.m_s_sync.d_data[40] ),
    .S(net204),
    .X(_1320_));
 sky130_fd_sc_hd__mux2_1 _1446_ (.A0(net601),
    .A1(\wb_cross_clk.m_s_sync.d_data[36] ),
    .S(_1313_),
    .X(_1321_));
 sky130_fd_sc_hd__or4_2 _1447_ (.A(_1318_),
    .B(_1319_),
    .C(_1320_),
    .D(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__mux2_1 _1448_ (.A0(net588),
    .A1(\wb_cross_clk.m_s_sync.d_data[41] ),
    .S(net204),
    .X(_1323_));
 sky130_fd_sc_hd__mux2_1 _1449_ (.A0(net606),
    .A1(\wb_cross_clk.m_s_sync.d_data[38] ),
    .S(net204),
    .X(_1324_));
 sky130_fd_sc_hd__mux2_1 _1450_ (.A0(_1259_),
    .A1(\wb_cross_clk.m_s_sync.d_data[35] ),
    .S(net568),
    .X(_1325_));
 sky130_fd_sc_hd__mux2_1 _1451_ (.A0(net631),
    .A1(\wb_cross_clk.m_s_sync.d_data[44] ),
    .S(_1313_),
    .X(_1326_));
 sky130_fd_sc_hd__or4_2 _1452_ (.A(_1323_),
    .B(_1324_),
    .C(net569),
    .D(_1326_),
    .X(_0368_));
 sky130_fd_sc_hd__o31ai_4 _1453_ (.A1(_1317_),
    .A2(_1322_),
    .A3(_0368_),
    .B1(_1289_),
    .Y(_0369_));
 sky130_fd_sc_hd__a211o_1 _1454_ (.A1(\wb_compressor.state[0] ),
    .A2(net638),
    .B1(net201),
    .C1(\wb_compressor.state[1] ),
    .X(_0010_));
 sky130_fd_sc_hd__buf_2 _1455_ (.A(net103),
    .X(_0370_));
 sky130_fd_sc_hd__xor2_1 _1456_ (.A(net894),
    .B(\wb_cross_clk.prev_xor_err ),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _1457_ (.A0(\wb_compressor.wb_err ),
    .A1(_0371_),
    .S(net204),
    .X(_0372_));
 sky130_fd_sc_hd__o21ai_1 _1458_ (.A1(net90),
    .A2(_0372_),
    .B1(_1270_),
    .Y(_0373_));
 sky130_fd_sc_hd__nand4b_4 _1459_ (.A_N(net90),
    .B(_1253_),
    .C(_1271_),
    .D(_1275_),
    .Y(_0374_));
 sky130_fd_sc_hd__or2_1 _1460_ (.A(_1262_),
    .B(_1267_),
    .X(_0375_));
 sky130_fd_sc_hd__or4b_1 _1461_ (.A(_1253_),
    .B(_1254_),
    .C(_1257_),
    .D_N(net90),
    .X(_0376_));
 sky130_fd_sc_hd__xnor2_1 _1462_ (.A(_1251_),
    .B(_1252_),
    .Y(_0377_));
 sky130_fd_sc_hd__or4_4 _1463_ (.A(_1250_),
    .B(_0375_),
    .C(_0376_),
    .D(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__nand2_4 _1464_ (.A(_0374_),
    .B(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__or3b_4 _1465_ (.A(_0373_),
    .B(_0379_),
    .C_N(_1280_),
    .X(_0380_));
 sky130_fd_sc_hd__buf_4 _1466_ (.A(_1270_),
    .X(_0381_));
 sky130_fd_sc_hd__nand3_1 _1467_ (.A(_0381_),
    .B(_1276_),
    .C(_1280_),
    .Y(_0382_));
 sky130_fd_sc_hd__inv_2 _1468_ (.A(_1285_),
    .Y(_0383_));
 sky130_fd_sc_hd__o2111ai_2 _1469_ (.A1(_1270_),
    .A2(_0383_),
    .B1(_0378_),
    .C1(_0374_),
    .D1(_1280_),
    .Y(_0384_));
 sky130_fd_sc_hd__a21o_1 _1470_ (.A1(_0374_),
    .A2(_0378_),
    .B1(iram_wb_ack),
    .X(_0385_));
 sky130_fd_sc_hd__xor2_1 _1471_ (.A(net891),
    .B(net907),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _1472_ (.A0(\wb_compressor.wb_ack ),
    .A1(_0386_),
    .S(net204),
    .X(_0387_));
 sky130_fd_sc_hd__and4_1 _1473_ (.A(_1270_),
    .B(_1276_),
    .C(_1280_),
    .D(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__a31oi_4 _1474_ (.A1(_0382_),
    .A2(_0384_),
    .A3(_0385_),
    .B1(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__or2b_1 _1475_ (.A(net878),
    .B_N(net862),
    .X(_0390_));
 sky130_fd_sc_hd__a211o_2 _1476_ (.A1(_0380_),
    .A2(_0389_),
    .B1(_1281_),
    .C1(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__nor2_1 _1477_ (.A(_0370_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__clkinv_4 _1478_ (.A(net103),
    .Y(_0393_));
 sky130_fd_sc_hd__buf_2 _1479_ (.A(\sspi.bit_cnt[3] ),
    .X(_0394_));
 sky130_fd_sc_hd__inv_2 _1480_ (.A(\sspi.bit_cnt[2] ),
    .Y(_0395_));
 sky130_fd_sc_hd__nand2_4 _1481_ (.A(net821),
    .B(net855),
    .Y(_0396_));
 sky130_fd_sc_hd__nor2_1 _1482_ (.A(_0395_),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__nand2_1 _1483_ (.A(_0394_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__or2_1 _1484_ (.A(net803),
    .B(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__or2_1 _1485_ (.A(_0390_),
    .B(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__nor2_1 _1486_ (.A(net782),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__a32o_1 _1487_ (.A1(_0393_),
    .A2(\sspi.state[5] ),
    .A3(_0390_),
    .B1(_0401_),
    .B2(net865),
    .X(_0402_));
 sky130_fd_sc_hd__a21o_1 _1488_ (.A1(net796),
    .A2(_0392_),
    .B1(net866),
    .X(_0007_));
 sky130_fd_sc_hd__nor2b_2 _1489_ (.A(\sspi.sy_clk[2] ),
    .B_N(net862),
    .Y(_0403_));
 sky130_fd_sc_hd__clkinv_2 _1490_ (.A(net92),
    .Y(_0404_));
 sky130_fd_sc_hd__nand2_1 _1491_ (.A(_0404_),
    .B(_0403_),
    .Y(_0405_));
 sky130_fd_sc_hd__clkbuf_4 _1492_ (.A(net103),
    .X(_0406_));
 sky130_fd_sc_hd__a221o_1 _1493_ (.A1(net869),
    .A2(_0403_),
    .B1(_0405_),
    .B2(net867),
    .C1(_0406_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_4 _1494_ (.A(_0393_),
    .X(_0407_));
 sky130_fd_sc_hd__a32o_1 _1495_ (.A1(_0407_),
    .A2(\sspi.state[7] ),
    .A3(_0400_),
    .B1(_0392_),
    .B2(net698),
    .X(_0009_));
 sky130_fd_sc_hd__buf_2 _1496_ (.A(net702),
    .X(_0408_));
 sky130_fd_sc_hd__a32o_1 _1497_ (.A1(net842),
    .A2(net92),
    .A3(_0403_),
    .B1(_0400_),
    .B2(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__and2_1 _1498_ (.A(_0407_),
    .B(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_1 _1499_ (.A(_0410_),
    .X(_0008_));
 sky130_fd_sc_hd__a32o_1 _1500_ (.A1(net796),
    .A2(_0407_),
    .A3(_0391_),
    .B1(_0401_),
    .B2(_0408_),
    .X(_0003_));
 sky130_fd_sc_hd__or2_2 _1501_ (.A(_0395_),
    .B(_0396_),
    .X(_0411_));
 sky130_fd_sc_hd__nor2_1 _1502_ (.A(_0394_),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__and3_1 _1503_ (.A(net803),
    .B(_0403_),
    .C(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__and2_1 _1504_ (.A(_0393_),
    .B(net826),
    .X(_0414_));
 sky130_fd_sc_hd__a32o_1 _1505_ (.A1(_0407_),
    .A2(net842),
    .A3(_0390_),
    .B1(_0413_),
    .B2(_0414_),
    .X(_0004_));
 sky130_fd_sc_hd__nand2_1 _1506_ (.A(_0393_),
    .B(\sspi.state[4] ),
    .Y(_0415_));
 sky130_fd_sc_hd__nor2_1 _1507_ (.A(_0406_),
    .B(_0405_),
    .Y(_0416_));
 sky130_fd_sc_hd__a2bb2o_1 _1508_ (.A1_N(_0413_),
    .A2_N(_0415_),
    .B1(_0416_),
    .B2(net867),
    .X(_0006_));
 sky130_fd_sc_hd__a32o_1 _1509_ (.A1(_0407_),
    .A2(net698),
    .A3(_0391_),
    .B1(_0416_),
    .B2(net842),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _1510_ (.A0(\m_arbiter.wb0_o_dat[8] ),
    .A1(net42),
    .S(_1225_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_2 _1511_ (.A(_0417_),
    .X(net145));
 sky130_fd_sc_hd__mux2_1 _1512_ (.A0(\m_arbiter.wb0_o_dat[9] ),
    .A1(net43),
    .S(_1225_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_2 _1513_ (.A(_0418_),
    .X(net146));
 sky130_fd_sc_hd__mux2_1 _1514_ (.A0(\m_arbiter.wb0_o_dat[10] ),
    .A1(net29),
    .S(_1225_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_2 _1515_ (.A(_0419_),
    .X(net132));
 sky130_fd_sc_hd__mux2_1 _1516_ (.A0(\m_arbiter.wb0_o_dat[11] ),
    .A1(net30),
    .S(_1229_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_2 _1517_ (.A(_0420_),
    .X(net133));
 sky130_fd_sc_hd__mux2_1 _1518_ (.A0(\m_arbiter.wb0_o_dat[12] ),
    .A1(net31),
    .S(_1229_),
    .X(_0421_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1519_ (.A(_0421_),
    .X(net134));
 sky130_fd_sc_hd__mux2_1 _1520_ (.A0(\m_arbiter.wb0_o_dat[13] ),
    .A1(net32),
    .S(_1229_),
    .X(_0422_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1521_ (.A(_0422_),
    .X(net135));
 sky130_fd_sc_hd__mux2_1 _1522_ (.A0(\m_arbiter.wb0_o_dat[14] ),
    .A1(net33),
    .S(_1229_),
    .X(_0423_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1523_ (.A(_0423_),
    .X(net136));
 sky130_fd_sc_hd__mux2_1 _1524_ (.A0(\m_arbiter.wb0_o_dat[15] ),
    .A1(net34),
    .S(_1229_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_2 _1525_ (.A(_0424_),
    .X(net137));
 sky130_fd_sc_hd__inv_2 _1526_ (.A(net126),
    .Y(_0425_));
 sky130_fd_sc_hd__or4_2 _1527_ (.A(_1245_),
    .B(_1250_),
    .C(_1255_),
    .D(_1278_),
    .X(_0426_));
 sky130_fd_sc_hd__nor4_4 _1528_ (.A(_0425_),
    .B(_1268_),
    .C(_1277_),
    .D(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__or3b_1 _1529_ (.A(net122),
    .B(_1269_),
    .C_N(net123),
    .X(_0428_));
 sky130_fd_sc_hd__nor3_4 _1530_ (.A(_1256_),
    .B(_1268_),
    .C(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__nor2_2 _1531_ (.A(_0427_),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__a22o_1 _1532_ (.A1(net172),
    .A2(_0427_),
    .B1(_0429_),
    .B2(net148),
    .X(_0431_));
 sky130_fd_sc_hd__a21oi_1 _1533_ (.A1(net66),
    .A2(_0430_),
    .B1(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__buf_6 _1534_ (.A(_1313_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _1535_ (.A0(\wb_compressor.wb_i_dat[0] ),
    .A1(\wb_cross_clk.m_wb_i_dat[0] ),
    .S(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__and3_1 _1536_ (.A(_0381_),
    .B(_1276_),
    .C(_1280_),
    .X(_0435_));
 sky130_fd_sc_hd__buf_2 _1537_ (.A(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_4 _1538_ (.A(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__a22oi_1 _1539_ (.A1(net48),
    .A2(_0379_),
    .B1(_0434_),
    .B2(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__o21ai_2 _1540_ (.A1(_0381_),
    .A2(_0432_),
    .B1(_0438_),
    .Y(net106));
 sky130_fd_sc_hd__a22o_1 _1541_ (.A1(net183),
    .A2(_0427_),
    .B1(_0430_),
    .B2(net77),
    .X(_0439_));
 sky130_fd_sc_hd__a21oi_1 _1542_ (.A1(net159),
    .A2(_0429_),
    .B1(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__buf_4 _1543_ (.A(_1313_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_2 _1544_ (.A0(\wb_compressor.wb_i_dat[1] ),
    .A1(\wb_cross_clk.m_wb_i_dat[1] ),
    .S(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__a22oi_1 _1545_ (.A1(net55),
    .A2(_0379_),
    .B1(_0442_),
    .B2(_0436_),
    .Y(_0443_));
 sky130_fd_sc_hd__o21ai_2 _1546_ (.A1(_0381_),
    .A2(_0440_),
    .B1(_0443_),
    .Y(net113));
 sky130_fd_sc_hd__a22o_1 _1547_ (.A1(net192),
    .A2(_0427_),
    .B1(_0430_),
    .B2(net86),
    .X(_0444_));
 sky130_fd_sc_hd__a21oi_1 _1548_ (.A1(net166),
    .A2(_0429_),
    .B1(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__mux2_2 _1549_ (.A0(\wb_compressor.wb_i_dat[2] ),
    .A1(\wb_cross_clk.m_wb_i_dat[2] ),
    .S(_0441_),
    .X(_0446_));
 sky130_fd_sc_hd__a22oi_1 _1550_ (.A1(net56),
    .A2(_0379_),
    .B1(_0446_),
    .B2(_0436_),
    .Y(_0447_));
 sky130_fd_sc_hd__o21ai_2 _1551_ (.A1(_0381_),
    .A2(_0445_),
    .B1(_0447_),
    .Y(net114));
 sky130_fd_sc_hd__a22o_1 _1552_ (.A1(net194),
    .A2(_0427_),
    .B1(_0430_),
    .B2(net93),
    .X(_0448_));
 sky130_fd_sc_hd__a21oi_1 _1553_ (.A1(net167),
    .A2(_0429_),
    .B1(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__mux2_1 _1554_ (.A0(\wb_compressor.wb_i_dat[3] ),
    .A1(\wb_cross_clk.m_wb_i_dat[3] ),
    .S(_0441_),
    .X(_0450_));
 sky130_fd_sc_hd__a22oi_1 _1555_ (.A1(net57),
    .A2(_0379_),
    .B1(_0450_),
    .B2(_0436_),
    .Y(_0451_));
 sky130_fd_sc_hd__o21ai_2 _1556_ (.A1(_0381_),
    .A2(_0449_),
    .B1(_0451_),
    .Y(net115));
 sky130_fd_sc_hd__a22o_1 _1557_ (.A1(net195),
    .A2(_0427_),
    .B1(_0429_),
    .B2(net168),
    .X(_0452_));
 sky130_fd_sc_hd__a21oi_1 _1558_ (.A1(net94),
    .A2(_0430_),
    .B1(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__mux2_1 _1559_ (.A0(\wb_compressor.wb_i_dat[4] ),
    .A1(\wb_cross_clk.m_wb_i_dat[4] ),
    .S(_0441_),
    .X(_0454_));
 sky130_fd_sc_hd__a22oi_1 _1560_ (.A1(net58),
    .A2(_0379_),
    .B1(_0454_),
    .B2(_0436_),
    .Y(_0455_));
 sky130_fd_sc_hd__o21ai_2 _1561_ (.A1(_0381_),
    .A2(_0453_),
    .B1(_0455_),
    .Y(net116));
 sky130_fd_sc_hd__a22o_1 _1562_ (.A1(net196),
    .A2(_0427_),
    .B1(_0429_),
    .B2(net169),
    .X(_0456_));
 sky130_fd_sc_hd__a21oi_1 _1563_ (.A1(net95),
    .A2(_0430_),
    .B1(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__mux2_1 _1564_ (.A0(\wb_compressor.wb_i_dat[5] ),
    .A1(\wb_cross_clk.m_wb_i_dat[5] ),
    .S(_0441_),
    .X(_0458_));
 sky130_fd_sc_hd__a22oi_1 _1565_ (.A1(net59),
    .A2(_0379_),
    .B1(_0458_),
    .B2(_0436_),
    .Y(_0459_));
 sky130_fd_sc_hd__o21ai_2 _1566_ (.A1(_0381_),
    .A2(_0457_),
    .B1(_0459_),
    .Y(net117));
 sky130_fd_sc_hd__a22o_1 _1567_ (.A1(net197),
    .A2(_0427_),
    .B1(_0429_),
    .B2(net170),
    .X(_0460_));
 sky130_fd_sc_hd__a21oi_2 _1568_ (.A1(net96),
    .A2(_0430_),
    .B1(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__mux2_2 _1569_ (.A0(\wb_compressor.wb_i_dat[6] ),
    .A1(\wb_cross_clk.m_wb_i_dat[6] ),
    .S(_0441_),
    .X(_0462_));
 sky130_fd_sc_hd__a22oi_2 _1570_ (.A1(net60),
    .A2(_0379_),
    .B1(_0462_),
    .B2(_0436_),
    .Y(_0463_));
 sky130_fd_sc_hd__o21ai_4 _1571_ (.A1(_0381_),
    .A2(_0461_),
    .B1(_0463_),
    .Y(net118));
 sky130_fd_sc_hd__a22o_1 _1572_ (.A1(net198),
    .A2(_0427_),
    .B1(_0429_),
    .B2(net171),
    .X(_0464_));
 sky130_fd_sc_hd__a21oi_2 _1573_ (.A1(net97),
    .A2(_0430_),
    .B1(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__mux2_2 _1574_ (.A0(\wb_compressor.wb_i_dat[7] ),
    .A1(\wb_cross_clk.m_wb_i_dat[7] ),
    .S(_0441_),
    .X(_0466_));
 sky130_fd_sc_hd__a22oi_2 _1575_ (.A1(net61),
    .A2(_0379_),
    .B1(_0466_),
    .B2(_0436_),
    .Y(_0467_));
 sky130_fd_sc_hd__o21ai_4 _1576_ (.A1(_0381_),
    .A2(_0465_),
    .B1(_0467_),
    .Y(net119));
 sky130_fd_sc_hd__buf_2 _1577_ (.A(_0379_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_8 _1578_ (.A(_0441_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_2 _1579_ (.A0(\wb_compressor.wb_i_dat[8] ),
    .A1(\wb_cross_clk.m_wb_i_dat[8] ),
    .S(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__a22o_1 _1580_ (.A1(net62),
    .A2(_0468_),
    .B1(_0470_),
    .B2(_0437_),
    .X(net120));
 sky130_fd_sc_hd__mux2_1 _1581_ (.A0(\wb_compressor.wb_i_dat[9] ),
    .A1(\wb_cross_clk.m_wb_i_dat[9] ),
    .S(_0469_),
    .X(_0471_));
 sky130_fd_sc_hd__a22o_1 _1582_ (.A1(net63),
    .A2(_0468_),
    .B1(_0471_),
    .B2(_0437_),
    .X(net121));
 sky130_fd_sc_hd__mux2_1 _1583_ (.A0(\wb_compressor.wb_i_dat[10] ),
    .A1(\wb_cross_clk.m_wb_i_dat[10] ),
    .S(_0469_),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _1584_ (.A1(net49),
    .A2(_0468_),
    .B1(_0472_),
    .B2(_0437_),
    .X(net107));
 sky130_fd_sc_hd__mux2_2 _1585_ (.A0(\wb_compressor.wb_i_dat[11] ),
    .A1(\wb_cross_clk.m_wb_i_dat[11] ),
    .S(_0433_),
    .X(_0473_));
 sky130_fd_sc_hd__a22o_1 _1586_ (.A1(net50),
    .A2(_0468_),
    .B1(_0473_),
    .B2(_0437_),
    .X(net108));
 sky130_fd_sc_hd__mux2_1 _1587_ (.A0(\wb_compressor.wb_i_dat[12] ),
    .A1(\wb_cross_clk.m_wb_i_dat[12] ),
    .S(_0433_),
    .X(_0474_));
 sky130_fd_sc_hd__a22o_1 _1588_ (.A1(net51),
    .A2(_0468_),
    .B1(_0474_),
    .B2(_0437_),
    .X(net109));
 sky130_fd_sc_hd__mux2_2 _1589_ (.A0(\wb_compressor.wb_i_dat[13] ),
    .A1(\wb_cross_clk.m_wb_i_dat[13] ),
    .S(_0433_),
    .X(_0475_));
 sky130_fd_sc_hd__a22o_1 _1590_ (.A1(net52),
    .A2(_0468_),
    .B1(_0475_),
    .B2(_0437_),
    .X(net110));
 sky130_fd_sc_hd__mux2_2 _1591_ (.A0(\wb_compressor.wb_i_dat[14] ),
    .A1(\wb_cross_clk.m_wb_i_dat[14] ),
    .S(_0433_),
    .X(_0476_));
 sky130_fd_sc_hd__a22o_1 _1592_ (.A1(net53),
    .A2(_0468_),
    .B1(_0476_),
    .B2(_0437_),
    .X(net111));
 sky130_fd_sc_hd__mux2_2 _1593_ (.A0(\wb_compressor.wb_i_dat[15] ),
    .A1(\wb_cross_clk.m_wb_i_dat[15] ),
    .S(_0433_),
    .X(_0477_));
 sky130_fd_sc_hd__a22o_1 _1594_ (.A1(net54),
    .A2(_0468_),
    .B1(_0477_),
    .B2(_0437_),
    .X(net112));
 sky130_fd_sc_hd__mux2_2 _1595_ (.A0(clknet_leaf_4_user_clock2),
    .A1(\clk_div.res_clk ),
    .S(\clk_div.clock_sel_r ),
    .X(_0478_));
 sky130_fd_sc_hd__buf_1 _1596_ (.A(_0478_),
    .X(net190));
 sky130_fd_sc_hd__mux2_4 _1597_ (.A0(net564),
    .A1(net47),
    .S(_1229_),
    .X(_0479_));
 sky130_fd_sc_hd__and3_2 _1598_ (.A(_1285_),
    .B(_0468_),
    .C(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_1 _1599_ (.A(_0480_),
    .X(net147));
 sky130_fd_sc_hd__o31a_1 _1600_ (.A1(_1317_),
    .A2(_1322_),
    .A3(_0368_),
    .B1(_1289_),
    .X(_0481_));
 sky130_fd_sc_hd__and3_1 _1601_ (.A(_1311_),
    .B(\wb_compressor.state[0] ),
    .C(net632),
    .X(_0482_));
 sky130_fd_sc_hd__clkbuf_1 _1602_ (.A(net633),
    .X(_0001_));
 sky130_fd_sc_hd__or2_1 _1603_ (.A(\wb_compressor.state[4] ),
    .B(\wb_compressor.state[5] ),
    .X(_0483_));
 sky130_fd_sc_hd__and3_1 _1604_ (.A(_1299_),
    .B(_1301_),
    .C(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__clkbuf_4 _1605_ (.A(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_4 _1606_ (.A(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__and2b_1 _1607_ (.A_N(_1296_),
    .B(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_1 _1608_ (.A(_0487_),
    .X(_0000_));
 sky130_fd_sc_hd__inv_2 _1609_ (.A(_1225_),
    .Y(_0488_));
 sky130_fd_sc_hd__nor2_1 _1610_ (.A(_0488_),
    .B(_0389_),
    .Y(net104));
 sky130_fd_sc_hd__nor2_1 _1611_ (.A(_0488_),
    .B(_0380_),
    .Y(net105));
 sky130_fd_sc_hd__nor2_1 _1612_ (.A(\wb_compressor.state[1] ),
    .B(net668),
    .Y(_0489_));
 sky130_fd_sc_hd__nor2_1 _1613_ (.A(\wb_compressor.state[4] ),
    .B(\wb_compressor.state[5] ),
    .Y(_0490_));
 sky130_fd_sc_hd__and2_1 _1614_ (.A(_0490_),
    .B(_0489_),
    .X(_0491_));
 sky130_fd_sc_hd__nor2_1 _1615_ (.A(net201),
    .B(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__o21a_1 _1616_ (.A1(net201),
    .A2(_0491_),
    .B1(net673),
    .X(_0493_));
 sky130_fd_sc_hd__a41o_1 _1617_ (.A1(net85),
    .A2(_1289_),
    .A3(_0489_),
    .A4(_0492_),
    .B1(_0493_),
    .X(_0019_));
 sky130_fd_sc_hd__xor2_1 _1618_ (.A(net917),
    .B(net933),
    .X(_0494_));
 sky130_fd_sc_hd__or2_1 _1619_ (.A(\wb_compressor.wb_ack ),
    .B(\wb_compressor.wb_err ),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_2 _1620_ (.A(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__buf_4 _1621_ (.A(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _1622_ (.A0(net856),
    .A1(_0494_),
    .S(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_1 _1623_ (.A(net857),
    .X(_0020_));
 sky130_fd_sc_hd__xor2_1 _1624_ (.A(net944),
    .B(\wb_compressor.wb_err ),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _1625_ (.A0(net744),
    .A1(_0499_),
    .S(_0497_),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_1 _1626_ (.A(net745),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _1627_ (.A0(net838),
    .A1(\wb_compressor.wb_i_dat[0] ),
    .S(_0497_),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_1 _1628_ (.A(net839),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _1629_ (.A0(net845),
    .A1(\wb_compressor.wb_i_dat[1] ),
    .S(_0497_),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_1 _1630_ (.A(net846),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _1631_ (.A0(net801),
    .A1(\wb_compressor.wb_i_dat[2] ),
    .S(_0497_),
    .X(_0503_));
 sky130_fd_sc_hd__clkbuf_1 _1632_ (.A(net802),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _1633_ (.A0(net819),
    .A1(\wb_compressor.wb_i_dat[3] ),
    .S(_0497_),
    .X(_0504_));
 sky130_fd_sc_hd__clkbuf_1 _1634_ (.A(net820),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _1635_ (.A0(net858),
    .A1(\wb_compressor.wb_i_dat[4] ),
    .S(_0497_),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_1 _1636_ (.A(net859),
    .X(_0026_));
 sky130_fd_sc_hd__buf_4 _1637_ (.A(_0496_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _1638_ (.A0(net748),
    .A1(\wb_compressor.wb_i_dat[5] ),
    .S(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_1 _1639_ (.A(net749),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _1640_ (.A0(net790),
    .A1(\wb_compressor.wb_i_dat[6] ),
    .S(_0506_),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_1 _1641_ (.A(net791),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _1642_ (.A0(net828),
    .A1(\wb_compressor.wb_i_dat[7] ),
    .S(_0506_),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_1 _1643_ (.A(net829),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _1644_ (.A0(net852),
    .A1(\wb_compressor.wb_i_dat[8] ),
    .S(_0506_),
    .X(_0510_));
 sky130_fd_sc_hd__clkbuf_1 _1645_ (.A(net853),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1646_ (.A0(net768),
    .A1(\wb_compressor.wb_i_dat[9] ),
    .S(_0506_),
    .X(_0511_));
 sky130_fd_sc_hd__clkbuf_1 _1647_ (.A(net769),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _1648_ (.A0(net739),
    .A1(\wb_compressor.wb_i_dat[10] ),
    .S(_0506_),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_1 _1649_ (.A(net740),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _1650_ (.A0(net814),
    .A1(\wb_compressor.wb_i_dat[11] ),
    .S(_0506_),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_1 _1651_ (.A(net815),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _1652_ (.A0(net760),
    .A1(\wb_compressor.wb_i_dat[12] ),
    .S(_0506_),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_1 _1653_ (.A(net761),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _1654_ (.A0(net840),
    .A1(\wb_compressor.wb_i_dat[13] ),
    .S(_0506_),
    .X(_0515_));
 sky130_fd_sc_hd__clkbuf_1 _1655_ (.A(net841),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _1656_ (.A0(net850),
    .A1(\wb_compressor.wb_i_dat[14] ),
    .S(_0506_),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_1 _1657_ (.A(net851),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _1658_ (.A0(net847),
    .A1(\wb_compressor.wb_i_dat[15] ),
    .S(_0496_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_1 _1659_ (.A(net848),
    .X(_0037_));
 sky130_fd_sc_hd__and3_1 _1660_ (.A(_1285_),
    .B(_0468_),
    .C(_0389_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _1661_ (.A(_0518_),
    .X(_0038_));
 sky130_fd_sc_hd__mux4_1 _1662_ (.A0(\clk_div.cnt[0] ),
    .A1(\clk_div.cnt[1] ),
    .A2(\clk_div.cnt[2] ),
    .A3(\clk_div.cnt[3] ),
    .S0(\clk_div.curr_div[0] ),
    .S1(\clk_div.curr_div[1] ),
    .X(_0519_));
 sky130_fd_sc_hd__mux4_1 _1663_ (.A0(\clk_div.cnt[4] ),
    .A1(\clk_div.cnt[5] ),
    .A2(\clk_div.cnt[6] ),
    .A3(\clk_div.cnt[7] ),
    .S0(\clk_div.curr_div[0] ),
    .S1(\clk_div.curr_div[1] ),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _1664_ (.A0(_0519_),
    .A1(_0520_),
    .S(\clk_div.curr_div[2] ),
    .X(_0521_));
 sky130_fd_sc_hd__inv_2 _1665_ (.A(\clk_div.curr_div[2] ),
    .Y(_0522_));
 sky130_fd_sc_hd__mux4_1 _1666_ (.A0(\clk_div.cnt[8] ),
    .A1(\clk_div.cnt[9] ),
    .A2(\clk_div.cnt[10] ),
    .A3(\clk_div.cnt[11] ),
    .S0(\clk_div.curr_div[0] ),
    .S1(\clk_div.curr_div[1] ),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _1667_ (.A0(\clk_div.cnt[12] ),
    .A1(\clk_div.cnt[13] ),
    .S(\clk_div.curr_div[0] ),
    .X(_0524_));
 sky130_fd_sc_hd__and2b_1 _1668_ (.A_N(\clk_div.curr_div[0] ),
    .B(\clk_div.cnt[14] ),
    .X(_0525_));
 sky130_fd_sc_hd__a21bo_1 _1669_ (.A1(\clk_div.curr_div[0] ),
    .A2(\clk_div.cnt[15] ),
    .B1_N(\clk_div.curr_div[1] ),
    .X(_0526_));
 sky130_fd_sc_hd__o221a_1 _1670_ (.A1(\clk_div.curr_div[1] ),
    .A2(_0524_),
    .B1(_0525_),
    .B2(_0526_),
    .C1(\clk_div.curr_div[2] ),
    .X(_0527_));
 sky130_fd_sc_hd__inv_2 _1671_ (.A(\clk_div.curr_div[3] ),
    .Y(_0528_));
 sky130_fd_sc_hd__a211o_1 _1672_ (.A1(_0522_),
    .A2(_0523_),
    .B1(_0527_),
    .C1(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__o21ai_4 _1673_ (.A1(\clk_div.curr_div[3] ),
    .A2(_0521_),
    .B1(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__buf_2 _1674_ (.A(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__xnor2_1 _1675_ (.A(net687),
    .B(_0531_),
    .Y(_0039_));
 sky130_fd_sc_hd__or2_1 _1676_ (.A(_1268_),
    .B(_1277_),
    .X(_0532_));
 sky130_fd_sc_hd__or3_1 _1677_ (.A(net126),
    .B(_0426_),
    .C(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__and3b_2 _1678_ (.A_N(_0533_),
    .B(_1284_),
    .C(_0479_),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _1679_ (.A0(net776),
    .A1(net131),
    .S(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_1 _1680_ (.A(_0535_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _1681_ (.A0(net843),
    .A1(net138),
    .S(_0534_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_1 _1682_ (.A(_0536_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _1683_ (.A0(net789),
    .A1(net139),
    .S(_0534_),
    .X(_0537_));
 sky130_fd_sc_hd__clkbuf_1 _1684_ (.A(_0537_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _1685_ (.A0(net816),
    .A1(net140),
    .S(_0534_),
    .X(_0538_));
 sky130_fd_sc_hd__clkbuf_1 _1686_ (.A(_0538_),
    .X(_0043_));
 sky130_fd_sc_hd__a21oi_1 _1687_ (.A1(net703),
    .A2(_0530_),
    .B1(_0534_),
    .Y(_0539_));
 sky130_fd_sc_hd__nor2_1 _1688_ (.A(_0406_),
    .B(net704),
    .Y(_0044_));
 sky130_fd_sc_hd__o211a_1 _1689_ (.A1(\clk_div.curr_div[3] ),
    .A2(_0521_),
    .B1(_0529_),
    .C1(\clk_div.next_div_val ),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _1690_ (.A0(net909),
    .A1(net776),
    .S(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__or2_1 _1691_ (.A(_0370_),
    .B(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__clkbuf_1 _1692_ (.A(_0542_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _1693_ (.A0(\clk_div.curr_div[1] ),
    .A1(net843),
    .S(_0540_),
    .X(_0543_));
 sky130_fd_sc_hd__and2_1 _1694_ (.A(_0407_),
    .B(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__clkbuf_1 _1695_ (.A(_0544_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _1696_ (.A0(net913),
    .A1(net789),
    .S(_0540_),
    .X(_0545_));
 sky130_fd_sc_hd__or2_1 _1697_ (.A(_0370_),
    .B(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__clkbuf_1 _1698_ (.A(_0546_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _1699_ (.A0(net932),
    .A1(net816),
    .S(_0540_),
    .X(_0547_));
 sky130_fd_sc_hd__and2_1 _1700_ (.A(_0407_),
    .B(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__clkbuf_1 _1701_ (.A(_0548_),
    .X(_0048_));
 sky130_fd_sc_hd__xor2_1 _1702_ (.A(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[2] ),
    .B(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ),
    .X(_0549_));
 sky130_fd_sc_hd__buf_4 _1703_ (.A(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__buf_4 _1704_ (.A(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _1705_ (.A0(\wb_cross_clk.m_s_sync.d_data[0] ),
    .A1(net516),
    .S(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__and2_1 _1706_ (.A(_1300_),
    .B(net517),
    .X(_0553_));
 sky130_fd_sc_hd__clkbuf_1 _1707_ (.A(net518),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _1708_ (.A0(\wb_cross_clk.m_s_sync.d_data[1] ),
    .A1(net441),
    .S(_0551_),
    .X(_0554_));
 sky130_fd_sc_hd__and2_1 _1709_ (.A(_1300_),
    .B(net442),
    .X(_0555_));
 sky130_fd_sc_hd__clkbuf_1 _1710_ (.A(net443),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _1711_ (.A0(\wb_cross_clk.m_s_sync.d_data[2] ),
    .A1(net534),
    .S(_0551_),
    .X(_0556_));
 sky130_fd_sc_hd__and2_1 _1712_ (.A(_1300_),
    .B(net535),
    .X(_0557_));
 sky130_fd_sc_hd__clkbuf_1 _1713_ (.A(net536),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _1714_ (.A0(\wb_cross_clk.m_s_sync.d_data[3] ),
    .A1(net504),
    .S(_0551_),
    .X(_0558_));
 sky130_fd_sc_hd__and2_1 _1715_ (.A(_1300_),
    .B(net505),
    .X(_0559_));
 sky130_fd_sc_hd__clkbuf_1 _1716_ (.A(net506),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1717_ (.A0(\wb_cross_clk.m_s_sync.d_data[4] ),
    .A1(net525),
    .S(_0551_),
    .X(_0560_));
 sky130_fd_sc_hd__and2_1 _1718_ (.A(_1300_),
    .B(net526),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_1 _1719_ (.A(net527),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _1720_ (.A0(\wb_cross_clk.m_s_sync.d_data[5] ),
    .A1(net453),
    .S(_0551_),
    .X(_0562_));
 sky130_fd_sc_hd__and2_1 _1721_ (.A(_1300_),
    .B(net454),
    .X(_0563_));
 sky130_fd_sc_hd__clkbuf_1 _1722_ (.A(net455),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _1723_ (.A0(\wb_cross_clk.m_s_sync.d_data[6] ),
    .A1(net489),
    .S(_0551_),
    .X(_0564_));
 sky130_fd_sc_hd__and2_1 _1724_ (.A(_1300_),
    .B(net490),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_1 _1725_ (.A(net491),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _1726_ (.A0(\wb_cross_clk.m_s_sync.d_data[7] ),
    .A1(net471),
    .S(_0551_),
    .X(_0566_));
 sky130_fd_sc_hd__and2_1 _1727_ (.A(_1300_),
    .B(net472),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_1 _1728_ (.A(net473),
    .X(_0056_));
 sky130_fd_sc_hd__buf_2 _1729_ (.A(_1299_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _1730_ (.A0(\wb_cross_clk.m_s_sync.d_data[8] ),
    .A1(net447),
    .S(_0551_),
    .X(_0569_));
 sky130_fd_sc_hd__and2_1 _1731_ (.A(_0568_),
    .B(net448),
    .X(_0570_));
 sky130_fd_sc_hd__clkbuf_1 _1732_ (.A(net449),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _1733_ (.A0(\wb_cross_clk.m_s_sync.d_data[9] ),
    .A1(net492),
    .S(_0551_),
    .X(_0571_));
 sky130_fd_sc_hd__and2_1 _1734_ (.A(_0568_),
    .B(net493),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_1 _1735_ (.A(net494),
    .X(_0058_));
 sky130_fd_sc_hd__buf_4 _1736_ (.A(_0550_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _1737_ (.A0(\wb_cross_clk.m_s_sync.d_data[10] ),
    .A1(net432),
    .S(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__and2_1 _1738_ (.A(_0568_),
    .B(net433),
    .X(_0575_));
 sky130_fd_sc_hd__clkbuf_1 _1739_ (.A(net434),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _1740_ (.A0(\wb_cross_clk.m_s_sync.d_data[11] ),
    .A1(net462),
    .S(_0573_),
    .X(_0576_));
 sky130_fd_sc_hd__and2_1 _1741_ (.A(_0568_),
    .B(net463),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_1 _1742_ (.A(net464),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1743_ (.A0(\wb_cross_clk.m_s_sync.d_data[12] ),
    .A1(net429),
    .S(_0573_),
    .X(_0578_));
 sky130_fd_sc_hd__and2_1 _1744_ (.A(_0568_),
    .B(net430),
    .X(_0579_));
 sky130_fd_sc_hd__clkbuf_1 _1745_ (.A(net431),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1746_ (.A0(\wb_cross_clk.m_s_sync.d_data[13] ),
    .A1(net468),
    .S(_0573_),
    .X(_0580_));
 sky130_fd_sc_hd__and2_1 _1747_ (.A(_0568_),
    .B(net469),
    .X(_0581_));
 sky130_fd_sc_hd__clkbuf_1 _1748_ (.A(net470),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1749_ (.A0(\wb_cross_clk.m_s_sync.d_data[14] ),
    .A1(net438),
    .S(_0573_),
    .X(_0582_));
 sky130_fd_sc_hd__and2_1 _1750_ (.A(_0568_),
    .B(net439),
    .X(_0583_));
 sky130_fd_sc_hd__clkbuf_1 _1751_ (.A(net440),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1752_ (.A0(\wb_cross_clk.m_s_sync.d_data[15] ),
    .A1(net507),
    .S(_0573_),
    .X(_0584_));
 sky130_fd_sc_hd__and2_1 _1753_ (.A(_0568_),
    .B(net508),
    .X(_0585_));
 sky130_fd_sc_hd__clkbuf_1 _1754_ (.A(net509),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1755_ (.A0(\wb_cross_clk.m_s_sync.d_data[16] ),
    .A1(net450),
    .S(_0573_),
    .X(_0586_));
 sky130_fd_sc_hd__and2_1 _1756_ (.A(_0568_),
    .B(net451),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_1 _1757_ (.A(net452),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1758_ (.A0(\wb_cross_clk.m_s_sync.d_data[17] ),
    .A1(net435),
    .S(_0573_),
    .X(_0588_));
 sky130_fd_sc_hd__and2_1 _1759_ (.A(_0568_),
    .B(net436),
    .X(_0589_));
 sky130_fd_sc_hd__clkbuf_1 _1760_ (.A(net437),
    .X(_0066_));
 sky130_fd_sc_hd__buf_2 _1761_ (.A(_1299_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _1762_ (.A0(\wb_cross_clk.m_s_sync.d_data[18] ),
    .A1(net474),
    .S(_0573_),
    .X(_0591_));
 sky130_fd_sc_hd__and2_1 _1763_ (.A(_0590_),
    .B(net475),
    .X(_0592_));
 sky130_fd_sc_hd__clkbuf_1 _1764_ (.A(net476),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1765_ (.A0(\wb_cross_clk.m_s_sync.d_data[19] ),
    .A1(net465),
    .S(_0573_),
    .X(_0593_));
 sky130_fd_sc_hd__and2_1 _1766_ (.A(_0590_),
    .B(net466),
    .X(_0594_));
 sky130_fd_sc_hd__clkbuf_1 _1767_ (.A(net467),
    .X(_0068_));
 sky130_fd_sc_hd__buf_4 _1768_ (.A(_0550_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _1769_ (.A0(\wb_cross_clk.m_s_sync.d_data[20] ),
    .A1(net495),
    .S(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__and2_1 _1770_ (.A(_0590_),
    .B(net496),
    .X(_0597_));
 sky130_fd_sc_hd__clkbuf_1 _1771_ (.A(net497),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1772_ (.A0(\wb_cross_clk.m_s_sync.d_data[21] ),
    .A1(net486),
    .S(_0595_),
    .X(_0598_));
 sky130_fd_sc_hd__and2_1 _1773_ (.A(_0590_),
    .B(net487),
    .X(_0599_));
 sky130_fd_sc_hd__clkbuf_1 _1774_ (.A(net488),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1775_ (.A0(\wb_cross_clk.m_s_sync.d_data[22] ),
    .A1(net537),
    .S(_0595_),
    .X(_0600_));
 sky130_fd_sc_hd__and2_1 _1776_ (.A(_0590_),
    .B(net538),
    .X(_0601_));
 sky130_fd_sc_hd__clkbuf_1 _1777_ (.A(net539),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1778_ (.A0(\wb_cross_clk.m_s_sync.d_data[23] ),
    .A1(net480),
    .S(_0595_),
    .X(_0602_));
 sky130_fd_sc_hd__and2_1 _1779_ (.A(_0590_),
    .B(net481),
    .X(_0603_));
 sky130_fd_sc_hd__clkbuf_1 _1780_ (.A(net482),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1781_ (.A0(\wb_cross_clk.m_s_sync.d_data[24] ),
    .A1(net498),
    .S(_0595_),
    .X(_0604_));
 sky130_fd_sc_hd__and2_1 _1782_ (.A(_0590_),
    .B(net499),
    .X(_0605_));
 sky130_fd_sc_hd__clkbuf_1 _1783_ (.A(net500),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1784_ (.A0(\wb_cross_clk.m_s_sync.d_data[25] ),
    .A1(net477),
    .S(_0595_),
    .X(_0606_));
 sky130_fd_sc_hd__and2_1 _1785_ (.A(_0590_),
    .B(net478),
    .X(_0607_));
 sky130_fd_sc_hd__clkbuf_1 _1786_ (.A(net479),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1787_ (.A0(\wb_cross_clk.m_s_sync.d_data[26] ),
    .A1(net444),
    .S(_0595_),
    .X(_0608_));
 sky130_fd_sc_hd__and2_1 _1788_ (.A(_0590_),
    .B(net445),
    .X(_0609_));
 sky130_fd_sc_hd__clkbuf_1 _1789_ (.A(net446),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _1790_ (.A0(\wb_cross_clk.m_s_sync.d_data[27] ),
    .A1(net426),
    .S(_0595_),
    .X(_0610_));
 sky130_fd_sc_hd__and2_1 _1791_ (.A(_0590_),
    .B(net427),
    .X(_0611_));
 sky130_fd_sc_hd__clkbuf_1 _1792_ (.A(net428),
    .X(_0076_));
 sky130_fd_sc_hd__buf_2 _1793_ (.A(_1299_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _1794_ (.A0(\wb_cross_clk.m_s_sync.d_data[28] ),
    .A1(net552),
    .S(_0595_),
    .X(_0613_));
 sky130_fd_sc_hd__and2_1 _1795_ (.A(_0612_),
    .B(net553),
    .X(_0614_));
 sky130_fd_sc_hd__clkbuf_1 _1796_ (.A(net554),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1797_ (.A0(\wb_cross_clk.m_s_sync.d_data[29] ),
    .A1(net531),
    .S(_0595_),
    .X(_0615_));
 sky130_fd_sc_hd__and2_1 _1798_ (.A(_0612_),
    .B(net532),
    .X(_0616_));
 sky130_fd_sc_hd__clkbuf_1 _1799_ (.A(net533),
    .X(_0078_));
 sky130_fd_sc_hd__buf_4 _1800_ (.A(_0549_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _1801_ (.A0(\wb_cross_clk.m_s_sync.d_data[30] ),
    .A1(net549),
    .S(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__and2_1 _1802_ (.A(_0612_),
    .B(net550),
    .X(_0619_));
 sky130_fd_sc_hd__clkbuf_1 _1803_ (.A(net551),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _1804_ (.A0(\wb_cross_clk.m_s_sync.d_data[31] ),
    .A1(net528),
    .S(_0617_),
    .X(_0620_));
 sky130_fd_sc_hd__and2_1 _1805_ (.A(_0612_),
    .B(net529),
    .X(_0621_));
 sky130_fd_sc_hd__clkbuf_1 _1806_ (.A(net530),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _1807_ (.A0(\wb_cross_clk.m_s_sync.d_data[32] ),
    .A1(net543),
    .S(_0617_),
    .X(_0622_));
 sky130_fd_sc_hd__and2_1 _1808_ (.A(_0612_),
    .B(net544),
    .X(_0623_));
 sky130_fd_sc_hd__clkbuf_1 _1809_ (.A(net545),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _1810_ (.A0(\wb_cross_clk.m_s_sync.d_data[33] ),
    .A1(net501),
    .S(_0617_),
    .X(_0624_));
 sky130_fd_sc_hd__and2_1 _1811_ (.A(_0612_),
    .B(net502),
    .X(_0625_));
 sky130_fd_sc_hd__clkbuf_1 _1812_ (.A(net503),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _1813_ (.A0(\wb_cross_clk.m_s_sync.d_data[34] ),
    .A1(net483),
    .S(_0617_),
    .X(_0626_));
 sky130_fd_sc_hd__and2_1 _1814_ (.A(_0612_),
    .B(net484),
    .X(_0627_));
 sky130_fd_sc_hd__clkbuf_1 _1815_ (.A(net485),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _1816_ (.A0(\wb_cross_clk.m_s_sync.d_data[35] ),
    .A1(net560),
    .S(_0617_),
    .X(_0628_));
 sky130_fd_sc_hd__and2_1 _1817_ (.A(_0612_),
    .B(net561),
    .X(_0629_));
 sky130_fd_sc_hd__clkbuf_1 _1818_ (.A(_0629_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _1819_ (.A0(\wb_cross_clk.m_s_sync.d_data[36] ),
    .A1(net562),
    .S(_0617_),
    .X(_0630_));
 sky130_fd_sc_hd__and2_1 _1820_ (.A(_0612_),
    .B(net563),
    .X(_0631_));
 sky130_fd_sc_hd__clkbuf_1 _1821_ (.A(_0631_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _1822_ (.A0(\wb_cross_clk.m_s_sync.d_data[37] ),
    .A1(net510),
    .S(_0617_),
    .X(_0632_));
 sky130_fd_sc_hd__and2_1 _1823_ (.A(_0612_),
    .B(net511),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_1 _1824_ (.A(net512),
    .X(_0086_));
 sky130_fd_sc_hd__buf_2 _1825_ (.A(_1299_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _1826_ (.A0(\wb_cross_clk.m_s_sync.d_data[38] ),
    .A1(net558),
    .S(_0617_),
    .X(_0635_));
 sky130_fd_sc_hd__and2_1 _1827_ (.A(_0634_),
    .B(net559),
    .X(_0636_));
 sky130_fd_sc_hd__clkbuf_1 _1828_ (.A(_0636_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _1829_ (.A0(\wb_cross_clk.m_s_sync.d_data[39] ),
    .A1(net546),
    .S(_0617_),
    .X(_0637_));
 sky130_fd_sc_hd__and2_1 _1830_ (.A(_0634_),
    .B(net547),
    .X(_0638_));
 sky130_fd_sc_hd__clkbuf_1 _1831_ (.A(net548),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _1832_ (.A0(\wb_cross_clk.m_s_sync.d_data[40] ),
    .A1(net513),
    .S(_0550_),
    .X(_0639_));
 sky130_fd_sc_hd__and2_1 _1833_ (.A(_0634_),
    .B(net514),
    .X(_0640_));
 sky130_fd_sc_hd__clkbuf_1 _1834_ (.A(net515),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1835_ (.A0(\wb_cross_clk.m_s_sync.d_data[41] ),
    .A1(net522),
    .S(_0550_),
    .X(_0641_));
 sky130_fd_sc_hd__and2_1 _1836_ (.A(_0634_),
    .B(net523),
    .X(_0642_));
 sky130_fd_sc_hd__clkbuf_1 _1837_ (.A(net524),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _1838_ (.A0(\wb_cross_clk.m_s_sync.d_data[42] ),
    .A1(net540),
    .S(_0550_),
    .X(_0643_));
 sky130_fd_sc_hd__and2_1 _1839_ (.A(_0634_),
    .B(net541),
    .X(_0644_));
 sky130_fd_sc_hd__clkbuf_1 _1840_ (.A(net542),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _1841_ (.A0(\wb_cross_clk.m_s_sync.d_data[43] ),
    .A1(net459),
    .S(_0550_),
    .X(_0645_));
 sky130_fd_sc_hd__and2_1 _1842_ (.A(_0634_),
    .B(net460),
    .X(_0646_));
 sky130_fd_sc_hd__clkbuf_1 _1843_ (.A(net461),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _1844_ (.A0(\wb_cross_clk.m_s_sync.d_data[44] ),
    .A1(net519),
    .S(_0550_),
    .X(_0647_));
 sky130_fd_sc_hd__and2_1 _1845_ (.A(_0634_),
    .B(net520),
    .X(_0648_));
 sky130_fd_sc_hd__clkbuf_1 _1846_ (.A(net521),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _1847_ (.A0(\wb_cross_clk.m_s_sync.d_data[45] ),
    .A1(net456),
    .S(_0550_),
    .X(_0649_));
 sky130_fd_sc_hd__and2_1 _1848_ (.A(_0634_),
    .B(net457),
    .X(_0650_));
 sky130_fd_sc_hd__clkbuf_1 _1849_ (.A(net458),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _1850_ (.A0(\wb_cross_clk.m_s_sync.d_data[46] ),
    .A1(net555),
    .S(_0550_),
    .X(_0651_));
 sky130_fd_sc_hd__and2_1 _1851_ (.A(_0634_),
    .B(net556),
    .X(_0652_));
 sky130_fd_sc_hd__clkbuf_1 _1852_ (.A(net557),
    .X(_0095_));
 sky130_fd_sc_hd__nor2_1 _1853_ (.A(_0371_),
    .B(_0386_),
    .Y(_0653_));
 sky130_fd_sc_hd__nor2_1 _1854_ (.A(_0406_),
    .B(net908),
    .Y(_0096_));
 sky130_fd_sc_hd__or3_1 _1855_ (.A(_1250_),
    .B(_1255_),
    .C(_1262_),
    .X(_0654_));
 sky130_fd_sc_hd__inv_2 _1856_ (.A(\wb_cross_clk.prev_ack ),
    .Y(_0655_));
 sky130_fd_sc_hd__or4_1 _1857_ (.A(\wb_cross_clk.m_burst_cnt[3] ),
    .B(\wb_cross_clk.m_burst_cnt[2] ),
    .C(\wb_cross_clk.m_burst_cnt[1] ),
    .D(\wb_cross_clk.m_burst_cnt[0] ),
    .X(_0656_));
 sky130_fd_sc_hd__a21oi_1 _1858_ (.A1(\wb_cross_clk.prev_stb ),
    .A2(_0655_),
    .B1(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__and4_1 _1859_ (.A(_0436_),
    .B(_1282_),
    .C(_0654_),
    .D(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_4 _1860_ (.A(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__a21oi_1 _1861_ (.A1(net423),
    .A2(_0659_),
    .B1(_0406_),
    .Y(_0660_));
 sky130_fd_sc_hd__o21a_1 _1862_ (.A1(net423),
    .A2(_0659_),
    .B1(_0660_),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _1863_ (.A(net423),
    .B(_1311_),
    .X(_0661_));
 sky130_fd_sc_hd__clkbuf_1 _1864_ (.A(net424),
    .X(_0098_));
 sky130_fd_sc_hd__and2_1 _1865_ (.A(_0634_),
    .B(net723),
    .X(_0662_));
 sky130_fd_sc_hd__clkbuf_1 _1866_ (.A(_0662_),
    .X(_0099_));
 sky130_fd_sc_hd__and2_1 _1867_ (.A(_1311_),
    .B(net883),
    .X(_0663_));
 sky130_fd_sc_hd__clkbuf_1 _1868_ (.A(_0663_),
    .X(_0100_));
 sky130_fd_sc_hd__buf_2 _1869_ (.A(_0393_),
    .X(_0664_));
 sky130_fd_sc_hd__xor2_4 _1870_ (.A(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[2] ),
    .B(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ),
    .X(_0665_));
 sky130_fd_sc_hd__buf_4 _1871_ (.A(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _1872_ (.A0(net891),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[0] ),
    .S(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__and2_1 _1873_ (.A(_0664_),
    .B(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__clkbuf_1 _1874_ (.A(_0668_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1875_ (.A0(net894),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[1] ),
    .S(_0666_),
    .X(_0669_));
 sky130_fd_sc_hd__and2_1 _1876_ (.A(_0664_),
    .B(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__clkbuf_1 _1877_ (.A(_0670_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _1878_ (.A0(net934),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[2] ),
    .S(_0666_),
    .X(_0671_));
 sky130_fd_sc_hd__and2_1 _1879_ (.A(_0664_),
    .B(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__clkbuf_1 _1880_ (.A(_0672_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1881_ (.A0(net928),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[3] ),
    .S(_0666_),
    .X(_0673_));
 sky130_fd_sc_hd__and2_1 _1882_ (.A(_0664_),
    .B(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_1 _1883_ (.A(_0674_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _1884_ (.A0(net922),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[4] ),
    .S(_0666_),
    .X(_0675_));
 sky130_fd_sc_hd__and2_1 _1885_ (.A(_0664_),
    .B(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__clkbuf_1 _1886_ (.A(_0676_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1887_ (.A0(net931),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[5] ),
    .S(_0666_),
    .X(_0677_));
 sky130_fd_sc_hd__and2_1 _1888_ (.A(_0664_),
    .B(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__clkbuf_1 _1889_ (.A(_0678_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _1890_ (.A0(net927),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[6] ),
    .S(_0666_),
    .X(_0679_));
 sky130_fd_sc_hd__and2_1 _1891_ (.A(_0664_),
    .B(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__clkbuf_1 _1892_ (.A(_0680_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1893_ (.A0(net925),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[7] ),
    .S(_0666_),
    .X(_0681_));
 sky130_fd_sc_hd__and2_1 _1894_ (.A(_0664_),
    .B(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__clkbuf_1 _1895_ (.A(_0682_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _1896_ (.A0(net935),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[8] ),
    .S(_0666_),
    .X(_0683_));
 sky130_fd_sc_hd__and2_1 _1897_ (.A(_0664_),
    .B(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__clkbuf_1 _1898_ (.A(_0684_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1899_ (.A0(net920),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[9] ),
    .S(_0666_),
    .X(_0685_));
 sky130_fd_sc_hd__and2_1 _1900_ (.A(_0664_),
    .B(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__clkbuf_1 _1901_ (.A(_0686_),
    .X(_0110_));
 sky130_fd_sc_hd__buf_2 _1902_ (.A(_0393_),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _1903_ (.A0(net919),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[10] ),
    .S(_0665_),
    .X(_0688_));
 sky130_fd_sc_hd__and2_1 _1904_ (.A(_0687_),
    .B(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__clkbuf_1 _1905_ (.A(_0689_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _1906_ (.A0(net937),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[11] ),
    .S(_0665_),
    .X(_0690_));
 sky130_fd_sc_hd__and2_1 _1907_ (.A(_0687_),
    .B(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__clkbuf_1 _1908_ (.A(_0691_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _1909_ (.A0(net929),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[12] ),
    .S(_0665_),
    .X(_0692_));
 sky130_fd_sc_hd__and2_1 _1910_ (.A(_0687_),
    .B(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__clkbuf_1 _1911_ (.A(_0693_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1912_ (.A0(net930),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[13] ),
    .S(_0665_),
    .X(_0694_));
 sky130_fd_sc_hd__and2_1 _1913_ (.A(_0687_),
    .B(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__clkbuf_1 _1914_ (.A(_0695_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _1915_ (.A0(net923),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[14] ),
    .S(_0665_),
    .X(_0696_));
 sky130_fd_sc_hd__and2_1 _1916_ (.A(_0687_),
    .B(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__clkbuf_1 _1917_ (.A(_0697_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _1918_ (.A0(net921),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[15] ),
    .S(_0665_),
    .X(_0698_));
 sky130_fd_sc_hd__and2_1 _1919_ (.A(_0687_),
    .B(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__clkbuf_1 _1920_ (.A(_0699_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _1921_ (.A0(net926),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[16] ),
    .S(_0665_),
    .X(_0700_));
 sky130_fd_sc_hd__and2_1 _1922_ (.A(_0687_),
    .B(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__clkbuf_1 _1923_ (.A(_0701_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _1924_ (.A0(net924),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[17] ),
    .S(_0665_),
    .X(_0702_));
 sky130_fd_sc_hd__and2_1 _1925_ (.A(_0687_),
    .B(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__clkbuf_1 _1926_ (.A(_0703_),
    .X(_0118_));
 sky130_fd_sc_hd__inv_2 _1927_ (.A(net757),
    .Y(_0704_));
 sky130_fd_sc_hd__mux2_1 _1928_ (.A0(net516),
    .A1(_0704_),
    .S(_0659_),
    .X(_0705_));
 sky130_fd_sc_hd__clkbuf_1 _1929_ (.A(_0705_),
    .X(_0119_));
 sky130_fd_sc_hd__and2_2 _1930_ (.A(_1229_),
    .B(net2),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _1931_ (.A0(net441),
    .A1(_0706_),
    .S(_0659_),
    .X(_0707_));
 sky130_fd_sc_hd__clkbuf_1 _1932_ (.A(_0707_),
    .X(_0120_));
 sky130_fd_sc_hd__and2_2 _1933_ (.A(_1225_),
    .B(net1),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _1934_ (.A0(net534),
    .A1(_0708_),
    .S(_0659_),
    .X(_0709_));
 sky130_fd_sc_hd__clkbuf_1 _1935_ (.A(_0709_),
    .X(_0121_));
 sky130_fd_sc_hd__or2_2 _1936_ (.A(_0488_),
    .B(net44),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _1937_ (.A0(net504),
    .A1(_0710_),
    .S(_0659_),
    .X(_0711_));
 sky130_fd_sc_hd__clkbuf_1 _1938_ (.A(_0711_),
    .X(_0122_));
 sky130_fd_sc_hd__or2_2 _1939_ (.A(_0488_),
    .B(net45),
    .X(_0712_));
 sky130_fd_sc_hd__buf_4 _1940_ (.A(_0658_),
    .X(_0713_));
 sky130_fd_sc_hd__buf_4 _1941_ (.A(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _1942_ (.A0(net525),
    .A1(_0712_),
    .S(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__clkbuf_1 _1943_ (.A(_0715_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1944_ (.A0(net453),
    .A1(_0479_),
    .S(_0714_),
    .X(_0716_));
 sky130_fd_sc_hd__clkbuf_1 _1945_ (.A(_0716_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _1946_ (.A0(net489),
    .A1(net131),
    .S(_0714_),
    .X(_0717_));
 sky130_fd_sc_hd__clkbuf_1 _1947_ (.A(_0717_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _1948_ (.A0(net471),
    .A1(net138),
    .S(_0714_),
    .X(_0718_));
 sky130_fd_sc_hd__clkbuf_1 _1949_ (.A(_0718_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1950_ (.A0(net447),
    .A1(net139),
    .S(_0714_),
    .X(_0719_));
 sky130_fd_sc_hd__clkbuf_1 _1951_ (.A(_0719_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _1952_ (.A0(net492),
    .A1(net140),
    .S(_0714_),
    .X(_0720_));
 sky130_fd_sc_hd__clkbuf_1 _1953_ (.A(_0720_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _1954_ (.A0(net432),
    .A1(net141),
    .S(_0714_),
    .X(_0721_));
 sky130_fd_sc_hd__clkbuf_1 _1955_ (.A(_0721_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _1956_ (.A0(net462),
    .A1(net142),
    .S(_0714_),
    .X(_0722_));
 sky130_fd_sc_hd__clkbuf_1 _1957_ (.A(_0722_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _1958_ (.A0(net429),
    .A1(net143),
    .S(_0714_),
    .X(_0723_));
 sky130_fd_sc_hd__clkbuf_1 _1959_ (.A(_0723_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _1960_ (.A0(net468),
    .A1(net144),
    .S(_0714_),
    .X(_0724_));
 sky130_fd_sc_hd__clkbuf_1 _1961_ (.A(_0724_),
    .X(_0132_));
 sky130_fd_sc_hd__buf_4 _1962_ (.A(_0713_),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _1963_ (.A0(net438),
    .A1(net145),
    .S(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__clkbuf_1 _1964_ (.A(_0726_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _1965_ (.A0(net507),
    .A1(net146),
    .S(_0725_),
    .X(_0727_));
 sky130_fd_sc_hd__clkbuf_1 _1966_ (.A(_0727_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _1967_ (.A0(net450),
    .A1(net132),
    .S(_0725_),
    .X(_0728_));
 sky130_fd_sc_hd__clkbuf_1 _1968_ (.A(_0728_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _1969_ (.A0(net435),
    .A1(net133),
    .S(_0725_),
    .X(_0729_));
 sky130_fd_sc_hd__clkbuf_1 _1970_ (.A(_0729_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _1971_ (.A0(net474),
    .A1(net134),
    .S(_0725_),
    .X(_0730_));
 sky130_fd_sc_hd__clkbuf_1 _1972_ (.A(_0730_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _1973_ (.A0(net465),
    .A1(net135),
    .S(_0725_),
    .X(_0731_));
 sky130_fd_sc_hd__clkbuf_1 _1974_ (.A(_0731_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _1975_ (.A0(net495),
    .A1(net136),
    .S(_0725_),
    .X(_0732_));
 sky130_fd_sc_hd__clkbuf_1 _1976_ (.A(_0732_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _1977_ (.A0(net486),
    .A1(net137),
    .S(_0725_),
    .X(_0733_));
 sky130_fd_sc_hd__clkbuf_1 _1978_ (.A(_0733_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _1979_ (.A0(net537),
    .A1(net122),
    .S(_0725_),
    .X(_0734_));
 sky130_fd_sc_hd__clkbuf_1 _1980_ (.A(_0734_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _1981_ (.A0(net480),
    .A1(net123),
    .S(_0725_),
    .X(_0735_));
 sky130_fd_sc_hd__clkbuf_1 _1982_ (.A(_0735_),
    .X(_0142_));
 sky130_fd_sc_hd__buf_4 _1983_ (.A(_0713_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _1984_ (.A0(net498),
    .A1(net124),
    .S(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__clkbuf_1 _1985_ (.A(_0737_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _1986_ (.A0(net477),
    .A1(net125),
    .S(_0736_),
    .X(_0738_));
 sky130_fd_sc_hd__clkbuf_1 _1987_ (.A(_0738_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _1988_ (.A0(net444),
    .A1(net126),
    .S(_0736_),
    .X(_0739_));
 sky130_fd_sc_hd__clkbuf_1 _1989_ (.A(_0739_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _1990_ (.A0(net426),
    .A1(net127),
    .S(_0736_),
    .X(_0740_));
 sky130_fd_sc_hd__clkbuf_1 _1991_ (.A(_0740_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _1992_ (.A0(net552),
    .A1(net128),
    .S(_0736_),
    .X(_0741_));
 sky130_fd_sc_hd__clkbuf_1 _1993_ (.A(_0741_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _1994_ (.A0(net531),
    .A1(net129),
    .S(_0736_),
    .X(_0742_));
 sky130_fd_sc_hd__clkbuf_1 _1995_ (.A(_0742_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _1996_ (.A0(net549),
    .A1(net812),
    .S(_0736_),
    .X(_0743_));
 sky130_fd_sc_hd__clkbuf_1 _1997_ (.A(_0743_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _1998_ (.A0(net528),
    .A1(_1265_),
    .S(_0736_),
    .X(_0744_));
 sky130_fd_sc_hd__clkbuf_1 _1999_ (.A(_0744_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2000_ (.A0(net543),
    .A1(_1264_),
    .S(_0736_),
    .X(_0745_));
 sky130_fd_sc_hd__clkbuf_1 _2001_ (.A(_0745_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2002_ (.A0(net501),
    .A1(_1266_),
    .S(_0736_),
    .X(_0746_));
 sky130_fd_sc_hd__clkbuf_1 _2003_ (.A(_0746_),
    .X(_0152_));
 sky130_fd_sc_hd__buf_4 _2004_ (.A(_0713_),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_1 _2005_ (.A0(net483),
    .A1(_1257_),
    .S(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__clkbuf_1 _2006_ (.A(_0748_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2007_ (.A0(net560),
    .A1(_1259_),
    .S(_0747_),
    .X(_0749_));
 sky130_fd_sc_hd__clkbuf_1 _2008_ (.A(_0749_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2009_ (.A0(net562),
    .A1(_1260_),
    .S(_0747_),
    .X(_0750_));
 sky130_fd_sc_hd__clkbuf_1 _2010_ (.A(_0750_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2011_ (.A0(net510),
    .A1(_1261_),
    .S(_0747_),
    .X(_0751_));
 sky130_fd_sc_hd__clkbuf_1 _2012_ (.A(_0751_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2013_ (.A0(net558),
    .A1(_1249_),
    .S(_0747_),
    .X(_0752_));
 sky130_fd_sc_hd__clkbuf_1 _2014_ (.A(_0752_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2015_ (.A0(net546),
    .A1(_1247_),
    .S(_0747_),
    .X(_0753_));
 sky130_fd_sc_hd__clkbuf_1 _2016_ (.A(_0753_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2017_ (.A0(net513),
    .A1(_1246_),
    .S(_0747_),
    .X(_0754_));
 sky130_fd_sc_hd__clkbuf_1 _2018_ (.A(_0754_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _2019_ (.A0(net522),
    .A1(_1248_),
    .S(_0747_),
    .X(_0755_));
 sky130_fd_sc_hd__clkbuf_1 _2020_ (.A(_0755_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2021_ (.A0(net540),
    .A1(_1252_),
    .S(_0747_),
    .X(_0756_));
 sky130_fd_sc_hd__clkbuf_1 _2022_ (.A(_0756_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2023_ (.A0(net459),
    .A1(_1253_),
    .S(_0747_),
    .X(_0757_));
 sky130_fd_sc_hd__clkbuf_1 _2024_ (.A(_0757_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2025_ (.A0(net519),
    .A1(_1254_),
    .S(_0713_),
    .X(_0758_));
 sky130_fd_sc_hd__clkbuf_1 _2026_ (.A(_0758_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2027_ (.A0(net456),
    .A1(_1251_),
    .S(_0713_),
    .X(_0759_));
 sky130_fd_sc_hd__clkbuf_1 _2028_ (.A(_0759_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2029_ (.A0(net555),
    .A1(_1284_),
    .S(_0713_),
    .X(_0760_));
 sky130_fd_sc_hd__clkbuf_1 _2030_ (.A(_0760_),
    .X(_0165_));
 sky130_fd_sc_hd__o21ai_1 _2031_ (.A1(net686),
    .A2(_0497_),
    .B1(_1300_),
    .Y(_0761_));
 sky130_fd_sc_hd__a21oi_1 _2032_ (.A1(net686),
    .A2(_0497_),
    .B1(_0761_),
    .Y(_0166_));
 sky130_fd_sc_hd__clkbuf_4 _2033_ (.A(_0393_),
    .X(_0762_));
 sky130_fd_sc_hd__and2_1 _2034_ (.A(\wb_cross_clk.s_m_sync.s_xfer_xor_flag ),
    .B(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__clkbuf_1 _2035_ (.A(_0763_),
    .X(_0167_));
 sky130_fd_sc_hd__and2_1 _2036_ (.A(_0687_),
    .B(net705),
    .X(_0764_));
 sky130_fd_sc_hd__clkbuf_1 _2037_ (.A(_0764_),
    .X(_0168_));
 sky130_fd_sc_hd__and2_1 _2038_ (.A(_0687_),
    .B(net916),
    .X(_0765_));
 sky130_fd_sc_hd__clkbuf_1 _2039_ (.A(_0765_),
    .X(_0169_));
 sky130_fd_sc_hd__and3_1 _2040_ (.A(_0762_),
    .B(_0437_),
    .C(_1282_),
    .X(_0766_));
 sky130_fd_sc_hd__clkbuf_1 _2041_ (.A(_0766_),
    .X(_0170_));
 sky130_fd_sc_hd__and2_1 _2042_ (.A(net894),
    .B(_0762_),
    .X(_0767_));
 sky130_fd_sc_hd__clkbuf_1 _2043_ (.A(_0767_),
    .X(_0171_));
 sky130_fd_sc_hd__xnor2_1 _2044_ (.A(net757),
    .B(_0659_),
    .Y(_0768_));
 sky130_fd_sc_hd__nor2_1 _2045_ (.A(_0406_),
    .B(_0768_),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _2046_ (.A(net565),
    .Y(_0769_));
 sky130_fd_sc_hd__nand3_1 _2047_ (.A(_0769_),
    .B(_0713_),
    .C(_0708_),
    .Y(_0770_));
 sky130_fd_sc_hd__nand3_1 _2048_ (.A(_0769_),
    .B(_0713_),
    .C(_0706_),
    .Y(_0771_));
 sky130_fd_sc_hd__xnor2_1 _2049_ (.A(\wb_cross_clk.m_burst_cnt[0] ),
    .B(_0653_),
    .Y(_0772_));
 sky130_fd_sc_hd__o21a_1 _2050_ (.A1(_0713_),
    .A2(_0772_),
    .B1(_0393_),
    .X(_0773_));
 sky130_fd_sc_hd__and3_1 _2051_ (.A(_0770_),
    .B(_0771_),
    .C(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__clkbuf_1 _2052_ (.A(_0774_),
    .X(_0173_));
 sky130_fd_sc_hd__or3_1 _2053_ (.A(\wb_cross_clk.m_burst_cnt[1] ),
    .B(net708),
    .C(_0653_),
    .X(_0775_));
 sky130_fd_sc_hd__o21ai_1 _2054_ (.A1(net708),
    .A2(_0653_),
    .B1(\wb_cross_clk.m_burst_cnt[1] ),
    .Y(_0776_));
 sky130_fd_sc_hd__a211oi_1 _2055_ (.A1(_0775_),
    .A2(net709),
    .B1(_0406_),
    .C1(_0659_),
    .Y(_0174_));
 sky130_fd_sc_hd__or2_1 _2056_ (.A(net892),
    .B(_0775_),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _2057_ (.A(net892),
    .B(_0775_),
    .Y(_0778_));
 sky130_fd_sc_hd__a211o_1 _2058_ (.A1(_0777_),
    .A2(_0778_),
    .B1(net103),
    .C1(_0659_),
    .X(_0779_));
 sky130_fd_sc_hd__o31ai_1 _2059_ (.A1(_0406_),
    .A2(_0706_),
    .A3(_0770_),
    .B1(_0779_),
    .Y(_0175_));
 sky130_fd_sc_hd__or2_1 _2060_ (.A(net885),
    .B(_0777_),
    .X(_0780_));
 sky130_fd_sc_hd__nand2_1 _2061_ (.A(net885),
    .B(_0777_),
    .Y(_0781_));
 sky130_fd_sc_hd__a21o_1 _2062_ (.A1(_0780_),
    .A2(_0781_),
    .B1(_0659_),
    .X(_0782_));
 sky130_fd_sc_hd__a21oi_1 _2063_ (.A1(_0771_),
    .A2(net886),
    .B1(_0406_),
    .Y(_0176_));
 sky130_fd_sc_hd__or3_1 _2064_ (.A(\wb_cross_clk.s_burst_cnt[2] ),
    .B(\wb_cross_clk.s_burst_cnt[1] ),
    .C(\wb_cross_clk.s_burst_cnt[0] ),
    .X(_0783_));
 sky130_fd_sc_hd__o21ai_1 _2065_ (.A1(\wb_cross_clk.s_burst_cnt[3] ),
    .A2(_0783_),
    .B1(_0496_),
    .Y(_0784_));
 sky130_fd_sc_hd__a21oi_1 _2066_ (.A1(\wb_cross_clk.m_s_sync.d_data[0] ),
    .A2(\wb_cross_clk.prev_xor_newreq ),
    .B1(_0496_),
    .Y(_0785_));
 sky130_fd_sc_hd__o21ai_1 _2067_ (.A1(\wb_cross_clk.m_s_sync.d_data[0] ),
    .A2(\wb_cross_clk.prev_xor_newreq ),
    .B1(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__and2_1 _2068_ (.A(_0784_),
    .B(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__nand2_1 _2069_ (.A(\wb_cross_clk.s_burst_cnt[0] ),
    .B(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__or2_1 _2070_ (.A(\wb_cross_clk.s_burst_cnt[0] ),
    .B(_0784_),
    .X(_0789_));
 sky130_fd_sc_hd__nor2_1 _2071_ (.A(\wb_cross_clk.m_s_sync.d_data[2] ),
    .B(\wb_cross_clk.m_s_sync.d_data[1] ),
    .Y(_0790_));
 sky130_fd_sc_hd__or3_1 _2072_ (.A(net565),
    .B(_0786_),
    .C(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__a31oi_1 _2073_ (.A1(_0788_),
    .A2(_0789_),
    .A3(net566),
    .B1(net201),
    .Y(_0177_));
 sky130_fd_sc_hd__and3_1 _2074_ (.A(net572),
    .B(_0786_),
    .C(_0789_),
    .X(_0792_));
 sky130_fd_sc_hd__o21ai_1 _2075_ (.A1(net572),
    .A2(_0789_),
    .B1(net566),
    .Y(_0793_));
 sky130_fd_sc_hd__o21a_1 _2076_ (.A1(_0792_),
    .A2(net573),
    .B1(_1312_),
    .X(_0178_));
 sky130_fd_sc_hd__inv_2 _2077_ (.A(_0787_),
    .Y(_0794_));
 sky130_fd_sc_hd__o21ai_1 _2078_ (.A1(net572),
    .A2(\wb_cross_clk.s_burst_cnt[0] ),
    .B1(net592),
    .Y(_0795_));
 sky130_fd_sc_hd__a21oi_1 _2079_ (.A1(_0783_),
    .A2(_0795_),
    .B1(_0784_),
    .Y(_0796_));
 sky130_fd_sc_hd__a31o_1 _2080_ (.A1(\wb_cross_clk.m_s_sync.d_data[1] ),
    .A2(_0769_),
    .A3(_0784_),
    .B1(_0787_),
    .X(_0797_));
 sky130_fd_sc_hd__buf_2 _2081_ (.A(_1311_),
    .X(_0798_));
 sky130_fd_sc_hd__o221a_1 _2082_ (.A1(net592),
    .A2(_0794_),
    .B1(_0796_),
    .B2(_0797_),
    .C1(_0798_),
    .X(_0179_));
 sky130_fd_sc_hd__a21o_1 _2083_ (.A1(_0496_),
    .A2(_0783_),
    .B1(_0787_),
    .X(_0799_));
 sky130_fd_sc_hd__and3_1 _2084_ (.A(net875),
    .B(_1311_),
    .C(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__clkbuf_1 _2085_ (.A(_0800_),
    .X(_0180_));
 sky130_fd_sc_hd__o211a_1 _2086_ (.A1(net884),
    .A2(_0497_),
    .B1(_0787_),
    .C1(_1312_),
    .X(_0181_));
 sky130_fd_sc_hd__and2_1 _2087_ (.A(_1311_),
    .B(net945),
    .X(_0801_));
 sky130_fd_sc_hd__clkbuf_1 _2088_ (.A(_0801_),
    .X(_0182_));
 sky130_fd_sc_hd__and2_1 _2089_ (.A(_1311_),
    .B(_0494_),
    .X(_0802_));
 sky130_fd_sc_hd__clkbuf_1 _2090_ (.A(_0802_),
    .X(_0183_));
 sky130_fd_sc_hd__and2_1 _2091_ (.A(net891),
    .B(_0762_),
    .X(_0803_));
 sky130_fd_sc_hd__clkbuf_1 _2092_ (.A(_0803_),
    .X(_0184_));
 sky130_fd_sc_hd__and2_1 _2093_ (.A(net872),
    .B(_1311_),
    .X(_0804_));
 sky130_fd_sc_hd__clkbuf_1 _2094_ (.A(_0804_),
    .X(_0185_));
 sky130_fd_sc_hd__buf_4 _2095_ (.A(_0441_),
    .X(_0805_));
 sky130_fd_sc_hd__mux2_1 _2096_ (.A0(net565),
    .A1(\wb_cross_clk.m_s_sync.d_data[5] ),
    .S(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__or2_1 _2097_ (.A(\wb_compressor.state[3] ),
    .B(\wb_compressor.state[6] ),
    .X(_0807_));
 sky130_fd_sc_hd__or2_2 _2098_ (.A(\wb_compressor.state[2] ),
    .B(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__or4_1 _2099_ (.A(net201),
    .B(\wb_compressor.state[1] ),
    .C(_0483_),
    .D(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__nor2_1 _2100_ (.A(net638),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__mux2_1 _2101_ (.A0(net575),
    .A1(_0806_),
    .S(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__clkbuf_1 _2102_ (.A(net576),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2103_ (.A0(_0708_),
    .A1(\wb_cross_clk.m_s_sync.d_data[2] ),
    .S(_0469_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_2 _2104_ (.A0(_0706_),
    .A1(\wb_cross_clk.m_s_sync.d_data[1] ),
    .S(_1313_),
    .X(_0813_));
 sky130_fd_sc_hd__or2_1 _2105_ (.A(_0812_),
    .B(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _2106_ (.A0(net676),
    .A1(_0814_),
    .S(_0810_),
    .X(_0815_));
 sky130_fd_sc_hd__clkbuf_1 _2107_ (.A(net677),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _2108_ (.A0(net666),
    .A1(_0813_),
    .S(_0810_),
    .X(_0816_));
 sky130_fd_sc_hd__clkbuf_1 _2109_ (.A(net667),
    .X(_0188_));
 sky130_fd_sc_hd__or3b_1 _2110_ (.A(_0490_),
    .B(_1290_),
    .C_N(_1296_),
    .X(_0817_));
 sky130_fd_sc_hd__nor2_1 _2111_ (.A(net915),
    .B(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__a2111o_1 _2112_ (.A1(_0369_),
    .A2(_0490_),
    .B1(_0808_),
    .C1(\wb_compressor.state[1] ),
    .D1(net201),
    .X(_0819_));
 sky130_fd_sc_hd__a21oi_1 _2113_ (.A1(_1290_),
    .A2(_0483_),
    .B1(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__mux2_1 _2114_ (.A0(net915),
    .A1(_0818_),
    .S(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__clkbuf_1 _2115_ (.A(_0821_),
    .X(_0189_));
 sky130_fd_sc_hd__and2_1 _2116_ (.A(\wb_compressor.burst_cnt[0] ),
    .B(\wb_compressor.burst_cnt[1] ),
    .X(_0822_));
 sky130_fd_sc_hd__nor3_1 _2117_ (.A(_1294_),
    .B(_0822_),
    .C(_0817_),
    .Y(_0823_));
 sky130_fd_sc_hd__mux2_1 _2118_ (.A0(net901),
    .A1(_0823_),
    .S(_0820_),
    .X(_0824_));
 sky130_fd_sc_hd__clkbuf_1 _2119_ (.A(_0824_),
    .X(_0190_));
 sky130_fd_sc_hd__o21a_1 _2120_ (.A1(_0822_),
    .A2(_0817_),
    .B1(net721),
    .X(_0825_));
 sky130_fd_sc_hd__nor3_1 _2121_ (.A(_1293_),
    .B(_0819_),
    .C(_0817_),
    .Y(_0826_));
 sky130_fd_sc_hd__o2bb2a_1 _2122_ (.A1_N(_0820_),
    .A2_N(_0825_),
    .B1(_0826_),
    .B2(net721),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _2123_ (.A0(net914),
    .A1(net67),
    .S(_0486_),
    .X(_0827_));
 sky130_fd_sc_hd__clkbuf_1 _2124_ (.A(_0827_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _2125_ (.A0(net904),
    .A1(net68),
    .S(_0486_),
    .X(_0828_));
 sky130_fd_sc_hd__clkbuf_1 _2126_ (.A(net905),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _2127_ (.A0(net897),
    .A1(net69),
    .S(_0486_),
    .X(_0829_));
 sky130_fd_sc_hd__clkbuf_1 _2128_ (.A(_0829_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _2129_ (.A0(net911),
    .A1(net70),
    .S(_0486_),
    .X(_0830_));
 sky130_fd_sc_hd__clkbuf_1 _2130_ (.A(net912),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _2131_ (.A0(net936),
    .A1(net71),
    .S(_0486_),
    .X(_0831_));
 sky130_fd_sc_hd__clkbuf_1 _2132_ (.A(_0831_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _2133_ (.A0(net900),
    .A1(net72),
    .S(_0486_),
    .X(_0832_));
 sky130_fd_sc_hd__clkbuf_1 _2134_ (.A(_0832_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _2135_ (.A0(net893),
    .A1(net73),
    .S(_0486_),
    .X(_0833_));
 sky130_fd_sc_hd__clkbuf_1 _2136_ (.A(_0833_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2137_ (.A0(net889),
    .A1(net74),
    .S(_0486_),
    .X(_0834_));
 sky130_fd_sc_hd__clkbuf_1 _2138_ (.A(_0834_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _2139_ (.A0(net895),
    .A1(net75),
    .S(_0485_),
    .X(_0835_));
 sky130_fd_sc_hd__clkbuf_1 _2140_ (.A(_0835_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2141_ (.A0(net902),
    .A1(net76),
    .S(_0485_),
    .X(_0836_));
 sky130_fd_sc_hd__clkbuf_1 _2142_ (.A(_0836_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2143_ (.A0(net910),
    .A1(net78),
    .S(_0485_),
    .X(_0837_));
 sky130_fd_sc_hd__clkbuf_1 _2144_ (.A(_0837_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _2145_ (.A0(net880),
    .A1(net79),
    .S(_0485_),
    .X(_0838_));
 sky130_fd_sc_hd__clkbuf_1 _2146_ (.A(_0838_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _2147_ (.A0(net906),
    .A1(net80),
    .S(_0485_),
    .X(_0839_));
 sky130_fd_sc_hd__clkbuf_1 _2148_ (.A(_0839_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _2149_ (.A0(net903),
    .A1(net81),
    .S(_0485_),
    .X(_0840_));
 sky130_fd_sc_hd__clkbuf_1 _2150_ (.A(_0840_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _2151_ (.A0(net898),
    .A1(net82),
    .S(_0485_),
    .X(_0841_));
 sky130_fd_sc_hd__clkbuf_1 _2152_ (.A(_0841_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _2153_ (.A0(net888),
    .A1(net83),
    .S(_0485_),
    .X(_0842_));
 sky130_fd_sc_hd__clkbuf_1 _2154_ (.A(_0842_),
    .X(_0207_));
 sky130_fd_sc_hd__and3_1 _2155_ (.A(net917),
    .B(_1299_),
    .C(_0491_),
    .X(_0843_));
 sky130_fd_sc_hd__a31o_1 _2156_ (.A1(net84),
    .A2(_0486_),
    .A3(_0489_),
    .B1(_0843_),
    .X(_0208_));
 sky130_fd_sc_hd__and2_1 _2157_ (.A(_0762_),
    .B(net91),
    .X(_0844_));
 sky130_fd_sc_hd__clkbuf_1 _2158_ (.A(_0844_),
    .X(_0209_));
 sky130_fd_sc_hd__and2_1 _2159_ (.A(_0762_),
    .B(net728),
    .X(_0845_));
 sky130_fd_sc_hd__clkbuf_1 _2160_ (.A(_0845_),
    .X(_0210_));
 sky130_fd_sc_hd__and2_1 _2161_ (.A(_0762_),
    .B(net862),
    .X(_0846_));
 sky130_fd_sc_hd__clkbuf_1 _2162_ (.A(_0846_),
    .X(_0211_));
 sky130_fd_sc_hd__inv_2 _2163_ (.A(\wb_compressor.state[1] ),
    .Y(_0847_));
 sky130_fd_sc_hd__a31o_1 _2164_ (.A1(_0847_),
    .A2(net638),
    .A3(_0490_),
    .B1(_0808_),
    .X(_0848_));
 sky130_fd_sc_hd__nand2_1 _2165_ (.A(net644),
    .B(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__or3_1 _2166_ (.A(net644),
    .B(_1290_),
    .C(_1296_),
    .X(_0850_));
 sky130_fd_sc_hd__a211o_1 _2167_ (.A1(_1297_),
    .A2(_0850_),
    .B1(_0808_),
    .C1(_0490_),
    .X(_0851_));
 sky130_fd_sc_hd__a21oi_1 _2168_ (.A1(net645),
    .A2(_0851_),
    .B1(net201),
    .Y(_0212_));
 sky130_fd_sc_hd__or2_2 _2169_ (.A(\wb_compressor.state[1] ),
    .B(\wb_compressor.state[4] ),
    .X(_0852_));
 sky130_fd_sc_hd__nor2_1 _2170_ (.A(\wb_compressor.state[2] ),
    .B(\wb_compressor.state[5] ),
    .Y(_0853_));
 sky130_fd_sc_hd__o211ai_1 _2171_ (.A1(_0852_),
    .A2(_0807_),
    .B1(_0853_),
    .C1(_1306_),
    .Y(_0854_));
 sky130_fd_sc_hd__nor2_4 _2172_ (.A(\wb_compressor.state[5] ),
    .B(_0808_),
    .Y(_0855_));
 sky130_fd_sc_hd__or3b_1 _2173_ (.A(net632),
    .B(_0852_),
    .C_N(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__a21o_1 _2174_ (.A1(_0853_),
    .A2(_0856_),
    .B1(net684),
    .X(_0857_));
 sky130_fd_sc_hd__and3_1 _2175_ (.A(_1311_),
    .B(_0854_),
    .C(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__clkbuf_1 _2176_ (.A(net685),
    .X(_0213_));
 sky130_fd_sc_hd__a211oi_4 _2177_ (.A1(_0369_),
    .A2(_0855_),
    .B1(_0852_),
    .C1(_1303_),
    .Y(_0859_));
 sky130_fd_sc_hd__buf_2 _2178_ (.A(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__buf_2 _2179_ (.A(_0855_),
    .X(_0861_));
 sky130_fd_sc_hd__a211o_2 _2180_ (.A1(_0369_),
    .A2(_0855_),
    .B1(_0852_),
    .C1(_1303_),
    .X(_0862_));
 sky130_fd_sc_hd__or3_4 _2181_ (.A(\wb_compressor.state[2] ),
    .B(\wb_compressor.state[5] ),
    .C(\wb_compressor.state[6] ),
    .X(_0863_));
 sky130_fd_sc_hd__mux2_1 _2182_ (.A0(net131),
    .A1(\wb_cross_clk.m_s_sync.d_data[6] ),
    .S(_0433_),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _2183_ (.A0(net122),
    .A1(\wb_cross_clk.m_s_sync.d_data[22] ),
    .S(_0433_),
    .X(_0865_));
 sky130_fd_sc_hd__a22o_1 _2184_ (.A1(_0863_),
    .A2(_0864_),
    .B1(net659),
    .B2(\wb_compressor.state[3] ),
    .X(_0866_));
 sky130_fd_sc_hd__or3_1 _2185_ (.A(_0861_),
    .B(_0862_),
    .C(net660),
    .X(_0867_));
 sky130_fd_sc_hd__o211a_1 _2186_ (.A1(net173),
    .A2(_0860_),
    .B1(net661),
    .C1(_1312_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _2187_ (.A0(net123),
    .A1(\wb_cross_clk.m_s_sync.d_data[23] ),
    .S(_0805_),
    .X(_0868_));
 sky130_fd_sc_hd__mux2_1 _2188_ (.A0(net138),
    .A1(\wb_cross_clk.m_s_sync.d_data[7] ),
    .S(_0433_),
    .X(_0869_));
 sky130_fd_sc_hd__buf_4 _2189_ (.A(_0441_),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_1 _2190_ (.A0(_0710_),
    .A1(\wb_cross_clk.m_s_sync.d_data[3] ),
    .S(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__a22o_1 _2191_ (.A1(_0863_),
    .A2(_0869_),
    .B1(_0871_),
    .B2(_0861_),
    .X(_0872_));
 sky130_fd_sc_hd__buf_2 _2192_ (.A(_0862_),
    .X(_0873_));
 sky130_fd_sc_hd__a211o_1 _2193_ (.A1(_1309_),
    .A2(net627),
    .B1(_0872_),
    .C1(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__o211a_1 _2194_ (.A1(net174),
    .A2(_0860_),
    .B1(net628),
    .C1(_1312_),
    .X(_0215_));
 sky130_fd_sc_hd__clkbuf_4 _2195_ (.A(_0863_),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _2196_ (.A0(net139),
    .A1(\wb_cross_clk.m_s_sync.d_data[8] ),
    .S(_0805_),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _2197_ (.A0(net124),
    .A1(\wb_cross_clk.m_s_sync.d_data[24] ),
    .S(_0433_),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _2198_ (.A0(_0712_),
    .A1(\wb_cross_clk.m_s_sync.d_data[4] ),
    .S(_0870_),
    .X(_0878_));
 sky130_fd_sc_hd__a22o_1 _2199_ (.A1(\wb_compressor.state[3] ),
    .A2(_0877_),
    .B1(_0878_),
    .B2(_0861_),
    .X(_0879_));
 sky130_fd_sc_hd__a211o_1 _2200_ (.A1(_0875_),
    .A2(net617),
    .B1(_0879_),
    .C1(_0873_),
    .X(_0880_));
 sky130_fd_sc_hd__o211a_1 _2201_ (.A1(net175),
    .A2(_0860_),
    .B1(net618),
    .C1(_1312_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _2202_ (.A0(net125),
    .A1(\wb_cross_clk.m_s_sync.d_data[25] ),
    .S(_0870_),
    .X(_0881_));
 sky130_fd_sc_hd__mux2_1 _2203_ (.A0(net140),
    .A1(\wb_cross_clk.m_s_sync.d_data[9] ),
    .S(_0805_),
    .X(_0882_));
 sky130_fd_sc_hd__a22o_1 _2204_ (.A1(_1309_),
    .A2(_0881_),
    .B1(net596),
    .B2(_0875_),
    .X(_0883_));
 sky130_fd_sc_hd__a211o_1 _2205_ (.A1(_0806_),
    .A2(_0861_),
    .B1(_0873_),
    .C1(net597),
    .X(_0884_));
 sky130_fd_sc_hd__o211a_1 _2206_ (.A1(net176),
    .A2(_0860_),
    .B1(net598),
    .C1(_1312_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2207_ (.A0(net126),
    .A1(\wb_cross_clk.m_s_sync.d_data[26] ),
    .S(_0469_),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _2208_ (.A0(net141),
    .A1(\wb_cross_clk.m_s_sync.d_data[10] ),
    .S(_0805_),
    .X(_0886_));
 sky130_fd_sc_hd__a22o_1 _2209_ (.A1(_1309_),
    .A2(_0885_),
    .B1(net653),
    .B2(_0875_),
    .X(_0887_));
 sky130_fd_sc_hd__a211o_1 _2210_ (.A1(_0813_),
    .A2(_0861_),
    .B1(_0873_),
    .C1(net654),
    .X(_0888_));
 sky130_fd_sc_hd__o211a_1 _2211_ (.A1(net177),
    .A2(_0860_),
    .B1(net655),
    .C1(_1312_),
    .X(_0218_));
 sky130_fd_sc_hd__inv_2 _2212_ (.A(_0813_),
    .Y(_0889_));
 sky130_fd_sc_hd__mux2_1 _2213_ (.A0(net127),
    .A1(\wb_cross_clk.m_s_sync.d_data[27] ),
    .S(_1313_),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _2214_ (.A0(net142),
    .A1(\wb_cross_clk.m_s_sync.d_data[11] ),
    .S(_1313_),
    .X(_0891_));
 sky130_fd_sc_hd__a22o_1 _2215_ (.A1(\wb_compressor.state[3] ),
    .A2(_0890_),
    .B1(net680),
    .B2(_0863_),
    .X(_0892_));
 sky130_fd_sc_hd__a31o_1 _2216_ (.A1(_0812_),
    .A2(_0889_),
    .A3(_0855_),
    .B1(net681),
    .X(_0893_));
 sky130_fd_sc_hd__or2_1 _2217_ (.A(_0862_),
    .B(net682),
    .X(_0894_));
 sky130_fd_sc_hd__o211a_1 _2218_ (.A1(net178),
    .A2(_0860_),
    .B1(_0894_),
    .C1(_1312_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _2219_ (.A0(net128),
    .A1(\wb_cross_clk.m_s_sync.d_data[28] ),
    .S(_0805_),
    .X(_0895_));
 sky130_fd_sc_hd__mux2_1 _2220_ (.A0(net143),
    .A1(\wb_cross_clk.m_s_sync.d_data[12] ),
    .S(_0805_),
    .X(_0896_));
 sky130_fd_sc_hd__a221o_1 _2221_ (.A1(_1309_),
    .A2(_0895_),
    .B1(net649),
    .B2(_0875_),
    .C1(_0862_),
    .X(_0897_));
 sky130_fd_sc_hd__o211a_1 _2222_ (.A1(net179),
    .A2(_0860_),
    .B1(net650),
    .C1(_1312_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _2223_ (.A0(net144),
    .A1(\wb_cross_clk.m_s_sync.d_data[13] ),
    .S(_0805_),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _2224_ (.A0(net129),
    .A1(\wb_cross_clk.m_s_sync.d_data[29] ),
    .S(_0805_),
    .X(_0899_));
 sky130_fd_sc_hd__a221o_1 _2225_ (.A1(_0875_),
    .A2(net641),
    .B1(_0899_),
    .B2(_1309_),
    .C1(_0862_),
    .X(_0900_));
 sky130_fd_sc_hd__o211a_1 _2226_ (.A1(net180),
    .A2(_0860_),
    .B1(net642),
    .C1(_0798_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _2227_ (.A0(_1263_),
    .A1(\wb_cross_clk.m_s_sync.d_data[30] ),
    .S(_0469_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _2228_ (.A0(net145),
    .A1(\wb_cross_clk.m_s_sync.d_data[14] ),
    .S(_0805_),
    .X(_0902_));
 sky130_fd_sc_hd__a22o_1 _2229_ (.A1(_1309_),
    .A2(_0901_),
    .B1(_0902_),
    .B2(_0875_),
    .X(_0903_));
 sky130_fd_sc_hd__a211o_1 _2230_ (.A1(net607),
    .A2(_0861_),
    .B1(_0873_),
    .C1(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__o211a_1 _2231_ (.A1(net181),
    .A2(_0860_),
    .B1(net608),
    .C1(_0798_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _2232_ (.A0(_1265_),
    .A1(\wb_cross_clk.m_s_sync.d_data[31] ),
    .S(_0469_),
    .X(_0905_));
 sky130_fd_sc_hd__mux2_1 _2233_ (.A0(net146),
    .A1(\wb_cross_clk.m_s_sync.d_data[15] ),
    .S(_0870_),
    .X(_0906_));
 sky130_fd_sc_hd__a22o_1 _2234_ (.A1(\wb_compressor.state[3] ),
    .A2(_0905_),
    .B1(_0906_),
    .B2(_0875_),
    .X(_0907_));
 sky130_fd_sc_hd__a211o_1 _2235_ (.A1(net622),
    .A2(_0861_),
    .B1(_0873_),
    .C1(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__o211a_1 _2236_ (.A1(net182),
    .A2(_0860_),
    .B1(net623),
    .C1(_0798_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _2237_ (.A0(_1264_),
    .A1(\wb_cross_clk.m_s_sync.d_data[32] ),
    .S(_0469_),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _2238_ (.A0(net132),
    .A1(\wb_cross_clk.m_s_sync.d_data[16] ),
    .S(_0870_),
    .X(_0910_));
 sky130_fd_sc_hd__a22o_1 _2239_ (.A1(\wb_compressor.state[3] ),
    .A2(_0909_),
    .B1(_0910_),
    .B2(_0863_),
    .X(_0911_));
 sky130_fd_sc_hd__a211o_1 _2240_ (.A1(net584),
    .A2(_0861_),
    .B1(_0873_),
    .C1(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__o211a_1 _2241_ (.A1(net184),
    .A2(_0859_),
    .B1(net585),
    .C1(_0798_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _2242_ (.A0(_1266_),
    .A1(\wb_cross_clk.m_s_sync.d_data[33] ),
    .S(_0469_),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _2243_ (.A0(net133),
    .A1(\wb_cross_clk.m_s_sync.d_data[17] ),
    .S(_0870_),
    .X(_0914_));
 sky130_fd_sc_hd__a22o_1 _2244_ (.A1(\wb_compressor.state[3] ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(_0863_),
    .X(_0915_));
 sky130_fd_sc_hd__a211o_1 _2245_ (.A1(net589),
    .A2(_0861_),
    .B1(_0873_),
    .C1(_0915_),
    .X(_0916_));
 sky130_fd_sc_hd__o211a_1 _2246_ (.A1(net185),
    .A2(_0859_),
    .B1(net590),
    .C1(_0798_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _2247_ (.A0(_1257_),
    .A1(\wb_cross_clk.m_s_sync.d_data[34] ),
    .S(_0469_),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _2248_ (.A0(net134),
    .A1(\wb_cross_clk.m_s_sync.d_data[18] ),
    .S(_0870_),
    .X(_0918_));
 sky130_fd_sc_hd__a22o_1 _2249_ (.A1(\wb_compressor.state[3] ),
    .A2(_0917_),
    .B1(_0918_),
    .B2(_0863_),
    .X(_0919_));
 sky130_fd_sc_hd__a211o_1 _2250_ (.A1(net612),
    .A2(_0861_),
    .B1(_0873_),
    .C1(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__o211a_1 _2251_ (.A1(net186),
    .A2(_0859_),
    .B1(net613),
    .C1(_0798_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _2252_ (.A0(net135),
    .A1(\wb_cross_clk.m_s_sync.d_data[19] ),
    .S(_0870_),
    .X(_0921_));
 sky130_fd_sc_hd__a22o_1 _2253_ (.A1(_1316_),
    .A2(_0855_),
    .B1(_0875_),
    .B2(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__a211o_1 _2254_ (.A1(_1309_),
    .A2(net569),
    .B1(_0873_),
    .C1(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__o211a_1 _2255_ (.A1(net187),
    .A2(_0859_),
    .B1(net570),
    .C1(_0798_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _2256_ (.A0(net136),
    .A1(\wb_cross_clk.m_s_sync.d_data[20] ),
    .S(_0870_),
    .X(_0924_));
 sky130_fd_sc_hd__a22o_1 _2257_ (.A1(_1326_),
    .A2(_0855_),
    .B1(_0875_),
    .B2(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__a211o_1 _2258_ (.A1(_1309_),
    .A2(net602),
    .B1(_0862_),
    .C1(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__o211a_1 _2259_ (.A1(net188),
    .A2(_0859_),
    .B1(net603),
    .C1(_0798_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _2260_ (.A0(net137),
    .A1(\wb_cross_clk.m_s_sync.d_data[21] ),
    .S(_0870_),
    .X(_0927_));
 sky130_fd_sc_hd__a22o_1 _2261_ (.A1(_1315_),
    .A2(_0855_),
    .B1(_0875_),
    .B2(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__a211o_1 _2262_ (.A1(_1309_),
    .A2(net579),
    .B1(_0862_),
    .C1(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__o211a_1 _2263_ (.A1(net189),
    .A2(_0859_),
    .B1(net580),
    .C1(_0798_),
    .X(_0229_));
 sky130_fd_sc_hd__a21o_2 _2264_ (.A1(_0380_),
    .A2(_0389_),
    .B1(_1281_),
    .X(_0930_));
 sky130_fd_sc_hd__inv_2 _2265_ (.A(\sspi.state[0] ),
    .Y(_0931_));
 sky130_fd_sc_hd__nand2_1 _2266_ (.A(_0931_),
    .B(_0403_),
    .Y(_0932_));
 sky130_fd_sc_hd__inv_2 _2267_ (.A(\sspi.state[5] ),
    .Y(_0933_));
 sky130_fd_sc_hd__a21oi_2 _2268_ (.A1(net698),
    .A2(_0933_),
    .B1(net796),
    .Y(_0934_));
 sky130_fd_sc_hd__or4_1 _2269_ (.A(\sspi.state[4] ),
    .B(\sspi.state[2] ),
    .C(\sspi.state[6] ),
    .D(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__nor2_1 _2270_ (.A(_0932_),
    .B(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__nand2_4 _2271_ (.A(_0393_),
    .B(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__buf_4 _2272_ (.A(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__o21ai_1 _2273_ (.A1(_0930_),
    .A2(_0938_),
    .B1(net688),
    .Y(_0939_));
 sky130_fd_sc_hd__or4_1 _2274_ (.A(_1225_),
    .B(_1281_),
    .C(_0380_),
    .D(_0937_),
    .X(_0940_));
 sky130_fd_sc_hd__nand2_1 _2275_ (.A(_0939_),
    .B(_0940_),
    .Y(_0230_));
 sky130_fd_sc_hd__a21oi_1 _2276_ (.A1(_0933_),
    .A2(\sspi.state[7] ),
    .B1(_0408_),
    .Y(_0941_));
 sky130_fd_sc_hd__a21oi_1 _2277_ (.A1(_0934_),
    .A2(_0941_),
    .B1(\sspi.state[2] ),
    .Y(_0942_));
 sky130_fd_sc_hd__o21bai_4 _2278_ (.A1(\sspi.state[4] ),
    .A2(_0942_),
    .B1_N(_0932_),
    .Y(_0943_));
 sky130_fd_sc_hd__nor2_1 _2279_ (.A(\sspi.state[1] ),
    .B(\sspi.state[3] ),
    .Y(_0944_));
 sky130_fd_sc_hd__nor3_2 _2280_ (.A(\sspi.state[4] ),
    .B(_0408_),
    .C(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__nor2_1 _2281_ (.A(_0943_),
    .B(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__inv_2 _2282_ (.A(net855),
    .Y(_0947_));
 sky130_fd_sc_hd__a211o_1 _2283_ (.A1(_0930_),
    .A2(_0945_),
    .B1(_0943_),
    .C1(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__clkbuf_4 _2284_ (.A(_0762_),
    .X(_0949_));
 sky130_fd_sc_hd__o211a_1 _2285_ (.A1(net855),
    .A2(_0946_),
    .B1(_0948_),
    .C1(_0949_),
    .X(_0231_));
 sky130_fd_sc_hd__or2_1 _2286_ (.A(_0943_),
    .B(_0945_),
    .X(_0950_));
 sky130_fd_sc_hd__o211a_1 _2287_ (.A1(_0930_),
    .A2(_0943_),
    .B1(_0950_),
    .C1(net821),
    .X(_0951_));
 sky130_fd_sc_hd__or2_2 _2288_ (.A(\sspi.bit_cnt[1] ),
    .B(\sspi.bit_cnt[0] ),
    .X(_0952_));
 sky130_fd_sc_hd__and3_1 _2289_ (.A(_0396_),
    .B(_0946_),
    .C(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__o21a_1 _2290_ (.A1(_0951_),
    .A2(_0953_),
    .B1(_0949_),
    .X(_0232_));
 sky130_fd_sc_hd__o211a_1 _2291_ (.A1(_0930_),
    .A2(_0943_),
    .B1(_0950_),
    .C1(net806),
    .X(_0954_));
 sky130_fd_sc_hd__or2_1 _2292_ (.A(_0396_),
    .B(_0943_),
    .X(_0955_));
 sky130_fd_sc_hd__a211oi_1 _2293_ (.A1(_0395_),
    .A2(_0955_),
    .B1(_0945_),
    .C1(_0397_),
    .Y(_0956_));
 sky130_fd_sc_hd__o21a_1 _2294_ (.A1(_0954_),
    .A2(_0956_),
    .B1(_0949_),
    .X(_0233_));
 sky130_fd_sc_hd__a31o_1 _2295_ (.A1(\sspi.bit_cnt[4] ),
    .A2(\sspi.state[4] ),
    .A3(_0412_),
    .B1(_0945_),
    .X(_0957_));
 sky130_fd_sc_hd__and2b_1 _2296_ (.A_N(_0957_),
    .B(_0398_),
    .X(_0958_));
 sky130_fd_sc_hd__a211o_1 _2297_ (.A1(_0930_),
    .A2(_0945_),
    .B1(_0958_),
    .C1(_0943_),
    .X(_0959_));
 sky130_fd_sc_hd__inv_2 _2298_ (.A(net783),
    .Y(_0960_));
 sky130_fd_sc_hd__o31ai_1 _2299_ (.A1(_0411_),
    .A2(_0943_),
    .A3(_0957_),
    .B1(_0960_),
    .Y(_0961_));
 sky130_fd_sc_hd__and3_1 _2300_ (.A(_0762_),
    .B(_0959_),
    .C(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__clkbuf_1 _2301_ (.A(_0962_),
    .X(_0234_));
 sky130_fd_sc_hd__or2_2 _2302_ (.A(\sspi.bit_cnt[2] ),
    .B(_0952_),
    .X(_0963_));
 sky130_fd_sc_hd__nor2_2 _2303_ (.A(net783),
    .B(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__and2_1 _2304_ (.A(net783),
    .B(_0963_),
    .X(_0965_));
 sky130_fd_sc_hd__or2_1 _2305_ (.A(_0964_),
    .B(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__buf_2 _2306_ (.A(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__nor2_1 _2307_ (.A(\sspi.state[4] ),
    .B(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__o22a_1 _2308_ (.A1(_0408_),
    .A2(_0944_),
    .B1(_0968_),
    .B2(_0411_),
    .X(_0969_));
 sky130_fd_sc_hd__a211o_1 _2309_ (.A1(_0930_),
    .A2(_0945_),
    .B1(_0969_),
    .C1(_0943_),
    .X(_0970_));
 sky130_fd_sc_hd__a2bb2o_1 _2310_ (.A1_N(_0399_),
    .A2_N(_0943_),
    .B1(net803),
    .B2(_0411_),
    .X(_0971_));
 sky130_fd_sc_hd__a32o_1 _2311_ (.A1(net803),
    .A2(_0407_),
    .A3(_0970_),
    .B1(_0971_),
    .B2(_0414_),
    .X(_0235_));
 sky130_fd_sc_hd__or3b_1 _2312_ (.A(net966),
    .B(\sspi.state[5] ),
    .C_N(net698),
    .X(_0972_));
 sky130_fd_sc_hd__clkinv_2 _2313_ (.A(\sspi.state[2] ),
    .Y(_0973_));
 sky130_fd_sc_hd__and4bb_1 _2314_ (.A_N(\sspi.state[4] ),
    .B_N(_0932_),
    .C(_0973_),
    .D(_0393_),
    .X(_0974_));
 sky130_fd_sc_hd__or3b_2 _2315_ (.A(_0972_),
    .B(_0408_),
    .C_N(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__nor3_4 _2316_ (.A(net103),
    .B(_0391_),
    .C(_0975_),
    .Y(_0976_));
 sky130_fd_sc_hd__clkbuf_4 _2317_ (.A(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__mux2_1 _2318_ (.A0(net879),
    .A1(net106),
    .S(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__clkbuf_1 _2319_ (.A(_0978_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _2320_ (.A0(net873),
    .A1(net113),
    .S(_0977_),
    .X(_0979_));
 sky130_fd_sc_hd__clkbuf_1 _2321_ (.A(_0979_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _2322_ (.A0(net877),
    .A1(net114),
    .S(_0977_),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_1 _2323_ (.A(_0980_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _2324_ (.A0(net876),
    .A1(net115),
    .S(_0977_),
    .X(_0981_));
 sky130_fd_sc_hd__clkbuf_1 _2325_ (.A(_0981_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _2326_ (.A0(net810),
    .A1(net116),
    .S(_0977_),
    .X(_0982_));
 sky130_fd_sc_hd__clkbuf_1 _2327_ (.A(_0982_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2328_ (.A0(net823),
    .A1(net117),
    .S(_0977_),
    .X(_0983_));
 sky130_fd_sc_hd__clkbuf_1 _2329_ (.A(_0983_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _2330_ (.A0(net837),
    .A1(net118),
    .S(_0977_),
    .X(_0984_));
 sky130_fd_sc_hd__clkbuf_1 _2331_ (.A(_0984_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _2332_ (.A0(net844),
    .A1(net119),
    .S(_0977_),
    .X(_0985_));
 sky130_fd_sc_hd__clkbuf_1 _2333_ (.A(_0985_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _2334_ (.A0(net780),
    .A1(net120),
    .S(_0977_),
    .X(_0986_));
 sky130_fd_sc_hd__clkbuf_1 _2335_ (.A(_0986_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _2336_ (.A0(net799),
    .A1(net121),
    .S(_0977_),
    .X(_0987_));
 sky130_fd_sc_hd__clkbuf_1 _2337_ (.A(_0987_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _2338_ (.A0(net860),
    .A1(net107),
    .S(_0976_),
    .X(_0988_));
 sky130_fd_sc_hd__clkbuf_1 _2339_ (.A(_0988_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _2340_ (.A0(net871),
    .A1(net108),
    .S(_0976_),
    .X(_0989_));
 sky130_fd_sc_hd__clkbuf_1 _2341_ (.A(_0989_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _2342_ (.A0(net887),
    .A1(net109),
    .S(_0976_),
    .X(_0990_));
 sky130_fd_sc_hd__clkbuf_1 _2343_ (.A(_0990_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _2344_ (.A0(net890),
    .A1(net110),
    .S(_0976_),
    .X(_0991_));
 sky130_fd_sc_hd__clkbuf_1 _2345_ (.A(_0991_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _2346_ (.A0(net899),
    .A1(net111),
    .S(_0976_),
    .X(_0992_));
 sky130_fd_sc_hd__clkbuf_1 _2347_ (.A(_0992_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _2348_ (.A0(net896),
    .A1(net112),
    .S(_0976_),
    .X(_0993_));
 sky130_fd_sc_hd__clkbuf_1 _2349_ (.A(_0993_),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_4 _2350_ (.A(net92),
    .X(_0994_));
 sky130_fd_sc_hd__and2_1 _2351_ (.A(_0408_),
    .B(_0974_),
    .X(_0995_));
 sky130_fd_sc_hd__buf_2 _2352_ (.A(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__nand2_1 _2353_ (.A(_0964_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__mux2_1 _2354_ (.A0(_0994_),
    .A1(net874),
    .S(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__clkbuf_1 _2355_ (.A(_0998_),
    .X(_0252_));
 sky130_fd_sc_hd__or2_2 _2356_ (.A(\sspi.bit_cnt[1] ),
    .B(_0947_),
    .X(_0999_));
 sky130_fd_sc_hd__or2_2 _2357_ (.A(\sspi.bit_cnt[2] ),
    .B(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__nand2_1 _2358_ (.A(_0408_),
    .B(_0974_),
    .Y(_1001_));
 sky130_fd_sc_hd__or2_2 _2359_ (.A(_0967_),
    .B(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__or2_1 _2360_ (.A(_1000_),
    .B(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__nor2_1 _2361_ (.A(_0404_),
    .B(_1000_),
    .Y(_1004_));
 sky130_fd_sc_hd__nor2_1 _2362_ (.A(_0967_),
    .B(_1001_),
    .Y(_1005_));
 sky130_fd_sc_hd__a22o_1 _2363_ (.A1(net720),
    .A2(_1003_),
    .B1(_1004_),
    .B2(_1005_),
    .X(_0253_));
 sky130_fd_sc_hd__nand2_2 _2364_ (.A(\sspi.bit_cnt[1] ),
    .B(_0947_),
    .Y(_1006_));
 sky130_fd_sc_hd__nor2_1 _2365_ (.A(net806),
    .B(net822),
    .Y(_1007_));
 sky130_fd_sc_hd__or2_2 _2366_ (.A(net835),
    .B(_1006_),
    .X(_1008_));
 sky130_fd_sc_hd__o21a_1 _2367_ (.A1(_1002_),
    .A2(_1008_),
    .B1(net742),
    .X(_1009_));
 sky130_fd_sc_hd__a31o_1 _2368_ (.A1(_0994_),
    .A2(_1005_),
    .A3(_1007_),
    .B1(_1009_),
    .X(_0254_));
 sky130_fd_sc_hd__or2_2 _2369_ (.A(\sspi.bit_cnt[2] ),
    .B(_0396_),
    .X(_1010_));
 sky130_fd_sc_hd__or2_1 _2370_ (.A(_1002_),
    .B(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__nor2_1 _2371_ (.A(_0404_),
    .B(_1010_),
    .Y(_1012_));
 sky130_fd_sc_hd__a22o_1 _2372_ (.A1(net724),
    .A2(_1011_),
    .B1(_1012_),
    .B2(_1005_),
    .X(_0255_));
 sky130_fd_sc_hd__nor2_1 _2373_ (.A(_0404_),
    .B(_0964_),
    .Y(_1013_));
 sky130_fd_sc_hd__or2_2 _2374_ (.A(_0395_),
    .B(_0952_),
    .X(_1014_));
 sky130_fd_sc_hd__nor2_1 _2375_ (.A(_1002_),
    .B(_1014_),
    .Y(_1015_));
 sky130_fd_sc_hd__mux2_1 _2376_ (.A0(net714),
    .A1(_1013_),
    .S(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__clkbuf_1 _2377_ (.A(_1016_),
    .X(_0256_));
 sky130_fd_sc_hd__buf_2 _2378_ (.A(_0394_),
    .X(_1017_));
 sky130_fd_sc_hd__or2_1 _2379_ (.A(_0395_),
    .B(_0999_),
    .X(_1018_));
 sky130_fd_sc_hd__nor2_1 _2380_ (.A(_1017_),
    .B(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__nand2_1 _2381_ (.A(_0996_),
    .B(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__mux2_1 _2382_ (.A0(_0994_),
    .A1(net797),
    .S(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__clkbuf_1 _2383_ (.A(_1021_),
    .X(_0257_));
 sky130_fd_sc_hd__or2_2 _2384_ (.A(_0395_),
    .B(_1006_),
    .X(_1022_));
 sky130_fd_sc_hd__nor2_1 _2385_ (.A(_1002_),
    .B(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__mux2_1 _2386_ (.A0(net813),
    .A1(_1013_),
    .S(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__clkbuf_1 _2387_ (.A(_1024_),
    .X(_0258_));
 sky130_fd_sc_hd__o21a_1 _2388_ (.A1(_0411_),
    .A2(_1002_),
    .B1(net770),
    .X(_1025_));
 sky130_fd_sc_hd__a31o_1 _2389_ (.A1(_0994_),
    .A2(_0397_),
    .A3(_1005_),
    .B1(_1025_),
    .X(_0259_));
 sky130_fd_sc_hd__nand2_2 _2390_ (.A(_0394_),
    .B(_0996_),
    .Y(_1026_));
 sky130_fd_sc_hd__or2_1 _2391_ (.A(_0963_),
    .B(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__mux2_1 _2392_ (.A0(_0994_),
    .A1(net817),
    .S(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__clkbuf_1 _2393_ (.A(_1028_),
    .X(_0260_));
 sky130_fd_sc_hd__o21a_1 _2394_ (.A1(_1000_),
    .A2(_1026_),
    .B1(net706),
    .X(_1029_));
 sky130_fd_sc_hd__a31o_1 _2395_ (.A1(_0967_),
    .A2(_0996_),
    .A3(_1004_),
    .B1(_1029_),
    .X(_0261_));
 sky130_fd_sc_hd__o21a_1 _2396_ (.A1(_1008_),
    .A2(_1026_),
    .B1(net827),
    .X(_1030_));
 sky130_fd_sc_hd__a41o_1 _2397_ (.A1(_0994_),
    .A2(_0965_),
    .A3(_0996_),
    .A4(_1007_),
    .B1(_1030_),
    .X(_0262_));
 sky130_fd_sc_hd__o21a_1 _2398_ (.A1(_1010_),
    .A2(_1026_),
    .B1(net794),
    .X(_1031_));
 sky130_fd_sc_hd__a31o_1 _2399_ (.A1(_0967_),
    .A2(_0996_),
    .A3(_1012_),
    .B1(_1031_),
    .X(_0263_));
 sky130_fd_sc_hd__or2_1 _2400_ (.A(_1014_),
    .B(_1026_),
    .X(_1032_));
 sky130_fd_sc_hd__nor4_1 _2401_ (.A(_0960_),
    .B(_0395_),
    .C(_0404_),
    .D(_0952_),
    .Y(_1033_));
 sky130_fd_sc_hd__a22o_1 _2402_ (.A1(net700),
    .A2(_1032_),
    .B1(_1033_),
    .B2(_0996_),
    .X(_0264_));
 sky130_fd_sc_hd__clkbuf_4 _2403_ (.A(net92),
    .X(_1034_));
 sky130_fd_sc_hd__or2_1 _2404_ (.A(_1018_),
    .B(_1026_),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _2405_ (.A0(_1034_),
    .A1(net773),
    .S(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__clkbuf_1 _2406_ (.A(_1036_),
    .X(_0265_));
 sky130_fd_sc_hd__or2_1 _2407_ (.A(_1022_),
    .B(_1026_),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _2408_ (.A0(_1034_),
    .A1(net785),
    .S(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__clkbuf_1 _2409_ (.A(_1038_),
    .X(_0266_));
 sky130_fd_sc_hd__or2_1 _2410_ (.A(_0398_),
    .B(_1001_),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(_1034_),
    .A1(net746),
    .S(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__clkbuf_1 _2412_ (.A(_1040_),
    .X(_0267_));
 sky130_fd_sc_hd__or2_1 _2413_ (.A(_0394_),
    .B(_0963_),
    .X(_1041_));
 sky130_fd_sc_hd__or2_1 _2414_ (.A(_0415_),
    .B(_0932_),
    .X(_1042_));
 sky130_fd_sc_hd__or3_1 _2415_ (.A(net803),
    .B(_1041_),
    .C(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__mux2_1 _2416_ (.A0(_1034_),
    .A1(net784),
    .S(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__clkbuf_1 _2417_ (.A(_1044_),
    .X(_0268_));
 sky130_fd_sc_hd__o21a_2 _2418_ (.A1(net807),
    .A2(_1041_),
    .B1(net92),
    .X(_1045_));
 sky130_fd_sc_hd__nor2_1 _2419_ (.A(_0415_),
    .B(_0932_),
    .Y(_1046_));
 sky130_fd_sc_hd__xnor2_1 _2420_ (.A(\sspi.bit_cnt[4] ),
    .B(_0964_),
    .Y(_1047_));
 sky130_fd_sc_hd__nand2_1 _2421_ (.A(_1046_),
    .B(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__or3_1 _2422_ (.A(_1017_),
    .B(_1000_),
    .C(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__mux2_1 _2423_ (.A0(_1045_),
    .A1(net788),
    .S(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__clkbuf_1 _2424_ (.A(_1050_),
    .X(_0269_));
 sky130_fd_sc_hd__or3_1 _2425_ (.A(_1017_),
    .B(_1008_),
    .C(_1048_),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_1 _2426_ (.A0(_1034_),
    .A1(net832),
    .S(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__clkbuf_1 _2427_ (.A(_1052_),
    .X(_0270_));
 sky130_fd_sc_hd__or3_1 _2428_ (.A(_1017_),
    .B(_1010_),
    .C(_1048_),
    .X(_1053_));
 sky130_fd_sc_hd__mux2_1 _2429_ (.A0(net804),
    .A1(net854),
    .S(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__clkbuf_1 _2430_ (.A(_1054_),
    .X(_0271_));
 sky130_fd_sc_hd__nor2_1 _2431_ (.A(_0394_),
    .B(_1014_),
    .Y(_1055_));
 sky130_fd_sc_hd__and3_1 _2432_ (.A(_1055_),
    .B(_1046_),
    .C(_1047_),
    .X(_1056_));
 sky130_fd_sc_hd__mux2_1 _2433_ (.A0(net743),
    .A1(net92),
    .S(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__clkbuf_1 _2434_ (.A(_1057_),
    .X(_0272_));
 sky130_fd_sc_hd__and2_1 _2435_ (.A(_1046_),
    .B(_1047_),
    .X(_1058_));
 sky130_fd_sc_hd__clkbuf_4 _2436_ (.A(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__nand2_1 _2437_ (.A(_1019_),
    .B(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(_1045_),
    .A1(net772),
    .S(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__clkbuf_1 _2439_ (.A(_1061_),
    .X(_0273_));
 sky130_fd_sc_hd__or3_1 _2440_ (.A(_1017_),
    .B(_1022_),
    .C(_1048_),
    .X(_1062_));
 sky130_fd_sc_hd__mux2_1 _2441_ (.A0(_1034_),
    .A1(net833),
    .S(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__clkbuf_1 _2442_ (.A(_1063_),
    .X(_0274_));
 sky130_fd_sc_hd__nand2_1 _2443_ (.A(_0412_),
    .B(_1059_),
    .Y(_1064_));
 sky130_fd_sc_hd__mux2_1 _2444_ (.A0(_1045_),
    .A1(net751),
    .S(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__clkbuf_1 _2445_ (.A(_1065_),
    .X(_0275_));
 sky130_fd_sc_hd__nand2_2 _2446_ (.A(_0394_),
    .B(_1059_),
    .Y(_1066_));
 sky130_fd_sc_hd__or2_1 _2447_ (.A(_0963_),
    .B(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__mux2_1 _2448_ (.A0(_1034_),
    .A1(net767),
    .S(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__clkbuf_1 _2449_ (.A(_1068_),
    .X(_0276_));
 sky130_fd_sc_hd__o21a_1 _2450_ (.A1(_1000_),
    .A2(_1066_),
    .B1(net733),
    .X(_1069_));
 sky130_fd_sc_hd__a31o_1 _2451_ (.A1(_0967_),
    .A2(_1004_),
    .A3(_1059_),
    .B1(_1069_),
    .X(_0277_));
 sky130_fd_sc_hd__o21a_1 _2452_ (.A1(_1008_),
    .A2(_1066_),
    .B1(net824),
    .X(_1070_));
 sky130_fd_sc_hd__a41o_1 _2453_ (.A1(_0994_),
    .A2(_0965_),
    .A3(_1007_),
    .A4(_1059_),
    .B1(_1070_),
    .X(_0278_));
 sky130_fd_sc_hd__o21a_1 _2454_ (.A1(_1010_),
    .A2(_1066_),
    .B1(net849),
    .X(_1071_));
 sky130_fd_sc_hd__a31o_1 _2455_ (.A1(_0967_),
    .A2(_1012_),
    .A3(_1059_),
    .B1(_1071_),
    .X(_0279_));
 sky130_fd_sc_hd__or2_1 _2456_ (.A(_1014_),
    .B(_1066_),
    .X(_1072_));
 sky130_fd_sc_hd__a22o_1 _2457_ (.A1(_1033_),
    .A2(_1059_),
    .B1(_1072_),
    .B2(net692),
    .X(_0280_));
 sky130_fd_sc_hd__or2_1 _2458_ (.A(_1018_),
    .B(_1066_),
    .X(_1073_));
 sky130_fd_sc_hd__mux2_1 _2459_ (.A0(_1034_),
    .A1(net763),
    .S(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__clkbuf_1 _2460_ (.A(_1074_),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _2461_ (.A(_1022_),
    .B(_1066_),
    .X(_1075_));
 sky130_fd_sc_hd__mux2_1 _2462_ (.A0(_1034_),
    .A1(net800),
    .S(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__clkbuf_1 _2463_ (.A(_1076_),
    .X(_0282_));
 sky130_fd_sc_hd__o21a_1 _2464_ (.A1(_0399_),
    .A2(_1042_),
    .B1(net758),
    .X(_1077_));
 sky130_fd_sc_hd__a41o_1 _2465_ (.A1(_1017_),
    .A2(_0994_),
    .A3(_0397_),
    .A4(_1059_),
    .B1(_1077_),
    .X(_0283_));
 sky130_fd_sc_hd__and3_1 _2466_ (.A(net807),
    .B(_0964_),
    .C(_1046_),
    .X(_1078_));
 sky130_fd_sc_hd__mux2_1 _2467_ (.A0(net805),
    .A1(net92),
    .S(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__clkbuf_1 _2468_ (.A(_1079_),
    .X(_0284_));
 sky130_fd_sc_hd__or2_2 _2469_ (.A(_1042_),
    .B(_1047_),
    .X(_1080_));
 sky130_fd_sc_hd__or3_1 _2470_ (.A(_1017_),
    .B(_1000_),
    .C(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__mux2_1 _2471_ (.A0(_1045_),
    .A1(net861),
    .S(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__clkbuf_1 _2472_ (.A(_1082_),
    .X(_0285_));
 sky130_fd_sc_hd__nor2_1 _2473_ (.A(_1042_),
    .B(_1047_),
    .Y(_1083_));
 sky130_fd_sc_hd__o31a_1 _2474_ (.A1(_1017_),
    .A2(_1008_),
    .A3(_1080_),
    .B1(net798),
    .X(_1084_));
 sky130_fd_sc_hd__a41o_1 _2475_ (.A1(_0960_),
    .A2(_0994_),
    .A3(_1007_),
    .A4(_1083_),
    .B1(_1084_),
    .X(_0286_));
 sky130_fd_sc_hd__or3_1 _2476_ (.A(_0394_),
    .B(_1010_),
    .C(_1080_),
    .X(_1085_));
 sky130_fd_sc_hd__mux2_1 _2477_ (.A0(_1045_),
    .A1(net792),
    .S(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__clkbuf_1 _2478_ (.A(_1086_),
    .X(_0287_));
 sky130_fd_sc_hd__o31a_1 _2479_ (.A1(_1017_),
    .A2(_1014_),
    .A3(_1080_),
    .B1(net868),
    .X(_1087_));
 sky130_fd_sc_hd__a31o_1 _2480_ (.A1(_0994_),
    .A2(_1055_),
    .A3(_1083_),
    .B1(_1087_),
    .X(_0288_));
 sky130_fd_sc_hd__o31a_1 _2481_ (.A1(_1017_),
    .A2(_1018_),
    .A3(_1080_),
    .B1(net716),
    .X(_1088_));
 sky130_fd_sc_hd__a31o_1 _2482_ (.A1(_1019_),
    .A2(net804),
    .A3(_1083_),
    .B1(_1088_),
    .X(_0289_));
 sky130_fd_sc_hd__or3_1 _2483_ (.A(_0394_),
    .B(_1022_),
    .C(_1080_),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_1 _2484_ (.A0(_1034_),
    .A1(net793),
    .S(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__clkbuf_1 _2485_ (.A(_1090_),
    .X(_0290_));
 sky130_fd_sc_hd__and3_1 _2486_ (.A(net803),
    .B(_0412_),
    .C(_1046_),
    .X(_1091_));
 sky130_fd_sc_hd__mux2_1 _2487_ (.A0(net825),
    .A1(_1013_),
    .S(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__clkbuf_1 _2488_ (.A(_1092_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _2489_ (.A0(net784),
    .A1(net657),
    .S(_0938_),
    .X(_1093_));
 sky130_fd_sc_hd__clkbuf_1 _2490_ (.A(_1093_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _2491_ (.A0(net788),
    .A1(net625),
    .S(_0938_),
    .X(_1094_));
 sky130_fd_sc_hd__clkbuf_1 _2492_ (.A(_1094_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _2493_ (.A0(net832),
    .A1(net781),
    .S(_0938_),
    .X(_1095_));
 sky130_fd_sc_hd__clkbuf_1 _2494_ (.A(_1095_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _2495_ (.A0(\sspi.req_addr[3] ),
    .A1(net808),
    .S(_0938_),
    .X(_1096_));
 sky130_fd_sc_hd__clkbuf_1 _2496_ (.A(net809),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _2497_ (.A0(net743),
    .A1(net765),
    .S(_0938_),
    .X(_1097_));
 sky130_fd_sc_hd__clkbuf_1 _2498_ (.A(_1097_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _2499_ (.A0(net772),
    .A1(net750),
    .S(_0938_),
    .X(_1098_));
 sky130_fd_sc_hd__clkbuf_1 _2500_ (.A(_1098_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _2501_ (.A0(net833),
    .A1(\m_arbiter.wb0_adr[6] ),
    .S(_0938_),
    .X(_1099_));
 sky130_fd_sc_hd__clkbuf_1 _2502_ (.A(net834),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _2503_ (.A0(net751),
    .A1(\m_arbiter.wb0_adr[7] ),
    .S(_0938_),
    .X(_1100_));
 sky130_fd_sc_hd__clkbuf_1 _2504_ (.A(net752),
    .X(_0299_));
 sky130_fd_sc_hd__buf_4 _2505_ (.A(_0937_),
    .X(_1101_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(net767),
    .A1(net811),
    .S(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__clkbuf_1 _2507_ (.A(_1102_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _2508_ (.A0(net733),
    .A1(\m_arbiter.wb0_adr[9] ),
    .S(_1101_),
    .X(_1103_));
 sky130_fd_sc_hd__clkbuf_1 _2509_ (.A(net734),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(net824),
    .A1(net818),
    .S(_1101_),
    .X(_1104_));
 sky130_fd_sc_hd__clkbuf_1 _2511_ (.A(_1104_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(net849),
    .A1(net741),
    .S(_1101_),
    .X(_1105_));
 sky130_fd_sc_hd__clkbuf_1 _2513_ (.A(_1105_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _2514_ (.A0(net692),
    .A1(net787),
    .S(_1101_),
    .X(_1106_));
 sky130_fd_sc_hd__clkbuf_1 _2515_ (.A(_1106_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _2516_ (.A0(net763),
    .A1(\m_arbiter.wb0_adr[13] ),
    .S(_1101_),
    .X(_1107_));
 sky130_fd_sc_hd__clkbuf_1 _2517_ (.A(net764),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _2518_ (.A0(net800),
    .A1(net600),
    .S(_1101_),
    .X(_1108_));
 sky130_fd_sc_hd__clkbuf_1 _2519_ (.A(_1108_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(net758),
    .A1(net577),
    .S(_1101_),
    .X(_1109_));
 sky130_fd_sc_hd__clkbuf_1 _2521_ (.A(_1109_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(net805),
    .A1(net605),
    .S(_1101_),
    .X(_1110_));
 sky130_fd_sc_hd__clkbuf_1 _2523_ (.A(_1110_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(net861),
    .A1(net620),
    .S(_1101_),
    .X(_1111_));
 sky130_fd_sc_hd__clkbuf_1 _2525_ (.A(_1111_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(net798),
    .A1(net582),
    .S(_0937_),
    .X(_1112_));
 sky130_fd_sc_hd__clkbuf_1 _2527_ (.A(_1112_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _2528_ (.A0(net792),
    .A1(net587),
    .S(_0937_),
    .X(_1113_));
 sky130_fd_sc_hd__clkbuf_1 _2529_ (.A(_1113_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(net868),
    .A1(net610),
    .S(_0937_),
    .X(_1114_));
 sky130_fd_sc_hd__clkbuf_1 _2531_ (.A(_1114_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2532_ (.A0(net716),
    .A1(net634),
    .S(_0937_),
    .X(_1115_));
 sky130_fd_sc_hd__clkbuf_1 _2533_ (.A(_1115_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2534_ (.A0(net793),
    .A1(net630),
    .S(_0937_),
    .X(_1116_));
 sky130_fd_sc_hd__clkbuf_1 _2535_ (.A(_1116_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _2536_ (.A0(net825),
    .A1(net771),
    .S(_0937_),
    .X(_1117_));
 sky130_fd_sc_hd__clkbuf_1 _2537_ (.A(_1117_),
    .X(_0315_));
 sky130_fd_sc_hd__inv_2 _2538_ (.A(_0938_),
    .Y(_1118_));
 sky130_fd_sc_hd__o21a_1 _2539_ (.A1(net564),
    .A2(_1118_),
    .B1(_0975_),
    .X(_0316_));
 sky130_fd_sc_hd__nand3b_4 _2540_ (.A_N(_0408_),
    .B(_0974_),
    .C(net796),
    .Y(_1119_));
 sky130_fd_sc_hd__buf_4 _2541_ (.A(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(net874),
    .A1(net775),
    .S(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__clkbuf_1 _2543_ (.A(_1121_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _2544_ (.A0(net720),
    .A1(net762),
    .S(_1120_),
    .X(_1122_));
 sky130_fd_sc_hd__clkbuf_1 _2545_ (.A(_1122_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(net742),
    .A1(net615),
    .S(_1120_),
    .X(_1123_));
 sky130_fd_sc_hd__clkbuf_1 _2547_ (.A(_1123_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(net724),
    .A1(net594),
    .S(_1120_),
    .X(_1124_));
 sky130_fd_sc_hd__clkbuf_1 _2549_ (.A(_1124_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(net714),
    .A1(net652),
    .S(_1120_),
    .X(_1125_));
 sky130_fd_sc_hd__clkbuf_1 _2551_ (.A(_1125_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _2552_ (.A0(net797),
    .A1(net678),
    .S(_1120_),
    .X(_1126_));
 sky130_fd_sc_hd__clkbuf_1 _2553_ (.A(_1126_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _2554_ (.A0(net813),
    .A1(net647),
    .S(_1120_),
    .X(_1127_));
 sky130_fd_sc_hd__clkbuf_1 _2555_ (.A(_1127_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _2556_ (.A0(net770),
    .A1(net640),
    .S(_1120_),
    .X(_1128_));
 sky130_fd_sc_hd__clkbuf_1 _2557_ (.A(_1128_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _2558_ (.A0(net817),
    .A1(net737),
    .S(_1120_),
    .X(_1129_));
 sky130_fd_sc_hd__clkbuf_1 _2559_ (.A(_1129_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _2560_ (.A0(net706),
    .A1(\m_arbiter.wb0_o_dat[9] ),
    .S(_1120_),
    .X(_1130_));
 sky130_fd_sc_hd__clkbuf_1 _2561_ (.A(net707),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _2562_ (.A0(\sspi.req_data[10] ),
    .A1(net778),
    .S(_1119_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_1 _2563_ (.A(net779),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _2564_ (.A0(net794),
    .A1(net759),
    .S(_1119_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _2565_ (.A(net795),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _2566_ (.A0(net700),
    .A1(net777),
    .S(_1119_),
    .X(_1133_));
 sky130_fd_sc_hd__clkbuf_1 _2567_ (.A(_1133_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _2568_ (.A0(net773),
    .A1(net766),
    .S(_1119_),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _2569_ (.A(net774),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _2570_ (.A0(net785),
    .A1(\m_arbiter.wb0_o_dat[14] ),
    .S(_1119_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_1 _2571_ (.A(net786),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(net746),
    .A1(\m_arbiter.wb0_o_dat[15] ),
    .S(_1119_),
    .X(_1136_));
 sky130_fd_sc_hd__clkbuf_1 _2573_ (.A(net747),
    .X(_0332_));
 sky130_fd_sc_hd__and2b_1 _2574_ (.A_N(net949),
    .B(_0530_),
    .X(_1137_));
 sky130_fd_sc_hd__clkbuf_1 _2575_ (.A(_1137_),
    .X(_0333_));
 sky130_fd_sc_hd__a21boi_1 _2576_ (.A1(\clk_div.cnt[0] ),
    .A2(net881),
    .B1_N(_0530_),
    .Y(_1138_));
 sky130_fd_sc_hd__o21a_1 _2577_ (.A1(\clk_div.cnt[0] ),
    .A2(net881),
    .B1(_1138_),
    .X(_0334_));
 sky130_fd_sc_hd__nand3_1 _2578_ (.A(\clk_div.cnt[0] ),
    .B(net881),
    .C(net940),
    .Y(_1139_));
 sky130_fd_sc_hd__a21o_1 _2579_ (.A1(\clk_div.cnt[0] ),
    .A2(\clk_div.cnt[1] ),
    .B1(net940),
    .X(_1140_));
 sky130_fd_sc_hd__and3_1 _2580_ (.A(_0530_),
    .B(net941),
    .C(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__clkbuf_1 _2581_ (.A(net942),
    .X(_0335_));
 sky130_fd_sc_hd__and4_1 _2582_ (.A(\clk_div.cnt[0] ),
    .B(\clk_div.cnt[1] ),
    .C(\clk_div.cnt[2] ),
    .D(\clk_div.cnt[3] ),
    .X(_1142_));
 sky130_fd_sc_hd__clkinv_2 _2583_ (.A(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__a31o_1 _2584_ (.A1(\clk_div.cnt[0] ),
    .A2(\clk_div.cnt[1] ),
    .A3(net940),
    .B1(net946),
    .X(_1144_));
 sky130_fd_sc_hd__and3_1 _2585_ (.A(_0530_),
    .B(_1143_),
    .C(net947),
    .X(_1145_));
 sky130_fd_sc_hd__clkbuf_1 _2586_ (.A(_1145_),
    .X(_0336_));
 sky130_fd_sc_hd__o21ai_1 _2587_ (.A1(net696),
    .A2(_1142_),
    .B1(_0531_),
    .Y(_1146_));
 sky130_fd_sc_hd__a21oi_1 _2588_ (.A1(net696),
    .A2(_1142_),
    .B1(_1146_),
    .Y(_0337_));
 sky130_fd_sc_hd__and3_1 _2589_ (.A(net696),
    .B(\clk_div.cnt[5] ),
    .C(_1142_),
    .X(_1147_));
 sky130_fd_sc_hd__clkinv_2 _2590_ (.A(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__a21o_1 _2591_ (.A1(net696),
    .A2(_1142_),
    .B1(net939),
    .X(_1149_));
 sky130_fd_sc_hd__and3_1 _2592_ (.A(_0530_),
    .B(_1148_),
    .C(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__clkbuf_1 _2593_ (.A(_1150_),
    .X(_0338_));
 sky130_fd_sc_hd__and2_1 _2594_ (.A(net755),
    .B(_1147_),
    .X(_1151_));
 sky130_fd_sc_hd__o21ai_1 _2595_ (.A1(net755),
    .A2(_1147_),
    .B1(_0531_),
    .Y(_1152_));
 sky130_fd_sc_hd__nor2_1 _2596_ (.A(_1151_),
    .B(net756),
    .Y(_0339_));
 sky130_fd_sc_hd__a21boi_1 _2597_ (.A1(net735),
    .A2(_1151_),
    .B1_N(_0530_),
    .Y(_1153_));
 sky130_fd_sc_hd__o21a_1 _2598_ (.A1(net735),
    .A2(_1151_),
    .B1(_1153_),
    .X(_0340_));
 sky130_fd_sc_hd__and3_1 _2599_ (.A(\clk_div.cnt[7] ),
    .B(\clk_div.cnt[8] ),
    .C(_1151_),
    .X(_1154_));
 sky130_fd_sc_hd__clkinv_2 _2600_ (.A(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__a31o_1 _2601_ (.A1(net755),
    .A2(net735),
    .A3(_1147_),
    .B1(net954),
    .X(_1156_));
 sky130_fd_sc_hd__and3_1 _2602_ (.A(_0530_),
    .B(_1155_),
    .C(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__clkbuf_1 _2603_ (.A(net955),
    .X(_0341_));
 sky130_fd_sc_hd__and2_1 _2604_ (.A(net729),
    .B(_1154_),
    .X(_1158_));
 sky130_fd_sc_hd__o21ai_1 _2605_ (.A1(net729),
    .A2(_1154_),
    .B1(_0531_),
    .Y(_1159_));
 sky130_fd_sc_hd__nor2_1 _2606_ (.A(_1158_),
    .B(net730),
    .Y(_0342_));
 sky130_fd_sc_hd__and3_1 _2607_ (.A(net729),
    .B(net717),
    .C(_1154_),
    .X(_1160_));
 sky130_fd_sc_hd__o21ai_1 _2608_ (.A1(net717),
    .A2(_1158_),
    .B1(_0531_),
    .Y(_1161_));
 sky130_fd_sc_hd__nor2_1 _2609_ (.A(_1160_),
    .B(net718),
    .Y(_0343_));
 sky130_fd_sc_hd__and2_1 _2610_ (.A(net732),
    .B(_1160_),
    .X(_1162_));
 sky130_fd_sc_hd__o21ai_1 _2611_ (.A1(net732),
    .A2(_1160_),
    .B1(_0531_),
    .Y(_1163_));
 sky130_fd_sc_hd__nor2_1 _2612_ (.A(_1162_),
    .B(_1163_),
    .Y(_0344_));
 sky130_fd_sc_hd__and3_1 _2613_ (.A(net732),
    .B(net711),
    .C(_1160_),
    .X(_1164_));
 sky130_fd_sc_hd__o21ai_1 _2614_ (.A1(net711),
    .A2(_1162_),
    .B1(_0531_),
    .Y(_1165_));
 sky130_fd_sc_hd__nor2_1 _2615_ (.A(_1164_),
    .B(net712),
    .Y(_0345_));
 sky130_fd_sc_hd__and2_1 _2616_ (.A(net738),
    .B(_1164_),
    .X(_1166_));
 sky130_fd_sc_hd__o21ai_1 _2617_ (.A1(net738),
    .A2(_1164_),
    .B1(_0531_),
    .Y(_1167_));
 sky130_fd_sc_hd__nor2_1 _2618_ (.A(_1166_),
    .B(_1167_),
    .Y(_0346_));
 sky130_fd_sc_hd__and3_1 _2619_ (.A(\clk_div.cnt[13] ),
    .B(net725),
    .C(_1164_),
    .X(_1168_));
 sky130_fd_sc_hd__o21ai_1 _2620_ (.A1(net725),
    .A2(_1166_),
    .B1(_0531_),
    .Y(_1169_));
 sky130_fd_sc_hd__nor2_1 _2621_ (.A(_1168_),
    .B(net726),
    .Y(_0347_));
 sky130_fd_sc_hd__o21a_1 _2622_ (.A1(net694),
    .A2(_1168_),
    .B1(_0531_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _2623_ (.A0(net715),
    .A1(_0930_),
    .S(_0936_),
    .X(_1170_));
 sky130_fd_sc_hd__and2_1 _2624_ (.A(_0762_),
    .B(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__clkbuf_1 _2625_ (.A(_1171_),
    .X(_0349_));
 sky130_fd_sc_hd__inv_2 _2626_ (.A(_0934_),
    .Y(_1172_));
 sky130_fd_sc_hd__or4_1 _2627_ (.A(\sspi.state[1] ),
    .B(\sspi.state[3] ),
    .C(\sspi.state[5] ),
    .D(\sspi.state[7] ),
    .X(_1173_));
 sky130_fd_sc_hd__or4b_1 _2628_ (.A(\sspi.state[4] ),
    .B(net842),
    .C(_0408_),
    .D_N(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__a21o_1 _2629_ (.A1(_0931_),
    .A2(_1174_),
    .B1(_0390_),
    .X(_1175_));
 sky130_fd_sc_hd__a21o_1 _2630_ (.A1(_0930_),
    .A2(_1172_),
    .B1(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__o221a_1 _2631_ (.A1(\sspi.res_data[6] ),
    .A2(_1006_),
    .B1(_0952_),
    .B2(\sspi.res_data[4] ),
    .C1(\sspi.bit_cnt[2] ),
    .X(_1177_));
 sky130_fd_sc_hd__o221a_1 _2632_ (.A1(\sspi.res_data[7] ),
    .A2(_0396_),
    .B1(_0999_),
    .B2(\sspi.res_data[5] ),
    .C1(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__o221a_1 _2633_ (.A1(\sspi.res_data[2] ),
    .A2(_1006_),
    .B1(_0952_),
    .B2(\sspi.res_data[0] ),
    .C1(_0395_),
    .X(_1179_));
 sky130_fd_sc_hd__o221a_1 _2634_ (.A1(\sspi.res_data[3] ),
    .A2(_0396_),
    .B1(_0999_),
    .B2(\sspi.res_data[1] ),
    .C1(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__or3_1 _2635_ (.A(_0394_),
    .B(_1178_),
    .C(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__o221a_1 _2636_ (.A1(\sspi.res_data[10] ),
    .A2(_1006_),
    .B1(_0952_),
    .B2(\sspi.res_data[8] ),
    .C1(_0395_),
    .X(_1182_));
 sky130_fd_sc_hd__o221a_1 _2637_ (.A1(\sspi.res_data[11] ),
    .A2(_0396_),
    .B1(_0999_),
    .B2(\sspi.res_data[9] ),
    .C1(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__o21a_1 _2638_ (.A1(\sspi.res_data[14] ),
    .A2(_1006_),
    .B1(\sspi.bit_cnt[2] ),
    .X(_1184_));
 sky130_fd_sc_hd__o22a_1 _2639_ (.A1(\sspi.res_data[15] ),
    .A2(_0396_),
    .B1(_0999_),
    .B2(\sspi.res_data[13] ),
    .X(_1185_));
 sky130_fd_sc_hd__o211a_1 _2640_ (.A1(\sspi.res_data[12] ),
    .A2(_0952_),
    .B1(_1184_),
    .C1(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__or3_1 _2641_ (.A(_0960_),
    .B(_1183_),
    .C(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__a21o_1 _2642_ (.A1(_1181_),
    .A2(_1187_),
    .B1(\sspi.state[5] ),
    .X(_1188_));
 sky130_fd_sc_hd__o211a_1 _2643_ (.A1(_0933_),
    .A2(net688),
    .B1(_0934_),
    .C1(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__o21ba_1 _2644_ (.A1(\sspi.state[0] ),
    .A2(_1189_),
    .B1_N(_1175_),
    .X(_1190_));
 sky130_fd_sc_hd__a211o_1 _2645_ (.A1(net863),
    .A2(_1176_),
    .B1(_1190_),
    .C1(_0406_),
    .X(_0350_));
 sky130_fd_sc_hd__nor4_1 _2646_ (.A(net122),
    .B(_1256_),
    .C(_1268_),
    .D(_1269_),
    .Y(_1191_));
 sky130_fd_sc_hd__and4_1 _2647_ (.A(net123),
    .B(_1285_),
    .C(_1191_),
    .D(_0479_),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_4 _2648_ (.A(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__mux2_1 _2649_ (.A0(net958),
    .A1(net131),
    .S(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__or2_1 _2650_ (.A(_0370_),
    .B(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__clkbuf_1 _2651_ (.A(_1195_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _2652_ (.A0(net960),
    .A1(net138),
    .S(_1193_),
    .X(_1196_));
 sky130_fd_sc_hd__or2_1 _2653_ (.A(_0370_),
    .B(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__clkbuf_1 _2654_ (.A(_1197_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _2655_ (.A0(net965),
    .A1(net139),
    .S(_1193_),
    .X(_1198_));
 sky130_fd_sc_hd__or2_1 _2656_ (.A(_0370_),
    .B(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__clkbuf_1 _2657_ (.A(_1199_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _2658_ (.A0(net963),
    .A1(net140),
    .S(_1193_),
    .X(_1200_));
 sky130_fd_sc_hd__or2_1 _2659_ (.A(_0370_),
    .B(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__clkbuf_1 _2660_ (.A(_1201_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _2661_ (.A0(net962),
    .A1(net141),
    .S(_1193_),
    .X(_1202_));
 sky130_fd_sc_hd__or2_1 _2662_ (.A(_0370_),
    .B(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__clkbuf_1 _2663_ (.A(_1203_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _2664_ (.A0(net959),
    .A1(net142),
    .S(_1193_),
    .X(_1204_));
 sky130_fd_sc_hd__or2_1 _2665_ (.A(_0370_),
    .B(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__clkbuf_1 _2666_ (.A(_1205_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _2667_ (.A0(net964),
    .A1(net143),
    .S(_1193_),
    .X(_1206_));
 sky130_fd_sc_hd__or2_1 _2668_ (.A(_0370_),
    .B(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__clkbuf_1 _2669_ (.A(_1207_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _2670_ (.A0(net961),
    .A1(net144),
    .S(_1193_),
    .X(_1208_));
 sky130_fd_sc_hd__or2_1 _2671_ (.A(net103),
    .B(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__clkbuf_1 _2672_ (.A(_1209_),
    .X(_0358_));
 sky130_fd_sc_hd__nand2_1 _2673_ (.A(_1285_),
    .B(_0479_),
    .Y(_1210_));
 sky130_fd_sc_hd__or4_1 _2674_ (.A(_0425_),
    .B(_0426_),
    .C(_0532_),
    .D(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__buf_2 _2675_ (.A(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__and3_2 _2676_ (.A(_1285_),
    .B(_0427_),
    .C(_0479_),
    .X(_1213_));
 sky130_fd_sc_hd__or2_1 _2677_ (.A(net951),
    .B(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__o211a_1 _2678_ (.A1(net131),
    .A2(_1212_),
    .B1(_1214_),
    .C1(_0949_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _2679_ (.A(net956),
    .B(_1213_),
    .X(_1215_));
 sky130_fd_sc_hd__o211a_1 _2680_ (.A1(net138),
    .A2(_1212_),
    .B1(_1215_),
    .C1(_0949_),
    .X(_0360_));
 sky130_fd_sc_hd__or2_1 _2681_ (.A(net953),
    .B(_1213_),
    .X(_1216_));
 sky130_fd_sc_hd__o211a_1 _2682_ (.A1(net139),
    .A2(_1212_),
    .B1(_1216_),
    .C1(_0949_),
    .X(_0361_));
 sky130_fd_sc_hd__or2_1 _2683_ (.A(net943),
    .B(_1213_),
    .X(_1217_));
 sky130_fd_sc_hd__o211a_1 _2684_ (.A1(net140),
    .A2(_1212_),
    .B1(_1217_),
    .C1(_0949_),
    .X(_0362_));
 sky130_fd_sc_hd__or2_1 _2685_ (.A(net952),
    .B(_1213_),
    .X(_1218_));
 sky130_fd_sc_hd__o211a_1 _2686_ (.A1(net141),
    .A2(_1212_),
    .B1(_1218_),
    .C1(_0949_),
    .X(_0363_));
 sky130_fd_sc_hd__or2_1 _2687_ (.A(net938),
    .B(_1213_),
    .X(_1219_));
 sky130_fd_sc_hd__o211a_1 _2688_ (.A1(net142),
    .A2(_1212_),
    .B1(_1219_),
    .C1(_0949_),
    .X(_0364_));
 sky130_fd_sc_hd__or2_1 _2689_ (.A(net950),
    .B(_1213_),
    .X(_1220_));
 sky130_fd_sc_hd__o211a_1 _2690_ (.A1(net143),
    .A2(_1212_),
    .B1(_1220_),
    .C1(_0949_),
    .X(_0365_));
 sky130_fd_sc_hd__or2_1 _2691_ (.A(net948),
    .B(_1213_),
    .X(_1221_));
 sky130_fd_sc_hd__o211a_1 _2692_ (.A1(net144),
    .A2(_1212_),
    .B1(_1221_),
    .C1(_0407_),
    .X(_0366_));
 sky130_fd_sc_hd__inv_2 _2693_ (.A(net65),
    .Y(_1222_));
 sky130_fd_sc_hd__a21oi_1 _2694_ (.A1(net64),
    .A2(_1222_),
    .B1(net98),
    .Y(_0015_));
 sky130_fd_sc_hd__a21oi_1 _2695_ (.A1(net64),
    .A2(_1222_),
    .B1(net98),
    .Y(_0016_));
 sky130_fd_sc_hd__a21oi_1 _2696_ (.A1(net64),
    .A2(_1222_),
    .B1(net98),
    .Y(_0017_));
 sky130_fd_sc_hd__a21oi_1 _2697_ (.A1(net64),
    .A2(_1222_),
    .B1(net98),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2_1 _2698_ (.A(net715),
    .B(_1283_),
    .Y(_1223_));
 sky130_fd_sc_hd__o211a_1 _2699_ (.A1(_1225_),
    .A2(net27),
    .B1(_0407_),
    .C1(_1223_),
    .X(_0367_));
 sky130_fd_sc_hd__dfxtp_1 _2700_ (.CLK(clknet_4_11_0_net190),
    .D(net674),
    .Q(\wb_compressor.wb_err ));
 sky130_fd_sc_hd__dfxtp_1 _2701_ (.CLK(clknet_leaf_4_user_clock2),
    .D(net90),
    .Q(\embed_s_ff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2702_ (.CLK(clknet_leaf_34_user_clock2),
    .D(net675),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _2703_ (.CLK(clknet_leaf_34_user_clock2),
    .D(net89),
    .Q(\disable_s_ff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2704_ (.CLK(clknet_leaf_34_user_clock2),
    .D(net664),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _2705_ (.CLK(clknet_leaf_11_user_clock2),
    .D(net88),
    .Q(\split_s_ff[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2706_ (.CLK(clknet_leaf_11_user_clock2),
    .D(net663),
    .Q(\clk_div.clock_sel ));
 sky130_fd_sc_hd__dfxtp_1 _2707_ (.CLK(clknet_leaf_34_user_clock2),
    .D(net87),
    .Q(\irq_s_ff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2708_ (.CLK(clknet_leaf_34_user_clock2),
    .D(net665),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_1 _2709_ (.CLK(clknet_4_9_0_net190),
    .D(_0020_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2710_ (.CLK(clknet_4_2_0_net190),
    .D(_0021_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2711_ (.CLK(clknet_4_10_0_net190),
    .D(_0022_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2712_ (.CLK(clknet_4_10_0_net190),
    .D(_0023_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2713_ (.CLK(clknet_4_10_0_net190),
    .D(_0024_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2714_ (.CLK(clknet_4_10_0_net190),
    .D(_0025_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2715_ (.CLK(clknet_4_8_0_net190),
    .D(_0026_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2716_ (.CLK(clknet_4_11_0_net190),
    .D(_0027_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2717_ (.CLK(clknet_4_11_0_net190),
    .D(_0028_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2718_ (.CLK(clknet_4_11_0_net190),
    .D(_0029_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2719_ (.CLK(clknet_4_14_0_net190),
    .D(_0030_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2720_ (.CLK(clknet_4_15_0_net190),
    .D(_0031_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2721_ (.CLK(clknet_4_13_0_net190),
    .D(_0032_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2722_ (.CLK(clknet_4_15_0_net190),
    .D(_0033_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2723_ (.CLK(clknet_4_13_0_net190),
    .D(_0034_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2724_ (.CLK(clknet_4_15_0_net190),
    .D(_0035_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2725_ (.CLK(clknet_4_15_0_net190),
    .D(_0036_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2726_ (.CLK(clknet_4_14_0_net190),
    .D(_0037_),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2727_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0038_),
    .Q(iram_wb_ack));
 sky130_fd_sc_hd__dfxtp_1 _2728_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0039_),
    .Q(\clk_div.res_clk ));
 sky130_fd_sc_hd__dfxtp_1 _2729_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0040_),
    .Q(\clk_div.next_div_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2730_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0041_),
    .Q(\clk_div.next_div_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2731_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0042_),
    .Q(\clk_div.next_div_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2732_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0043_),
    .Q(\clk_div.next_div_buff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2733_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0044_),
    .Q(\clk_div.next_div_val ));
 sky130_fd_sc_hd__dfxtp_2 _2734_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0045_),
    .Q(\clk_div.curr_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2735_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0046_),
    .Q(\clk_div.curr_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2736_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0047_),
    .Q(\clk_div.curr_div[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2737_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0048_),
    .Q(\clk_div.curr_div[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2738_ (.CLK(clknet_leaf_3_user_clock2),
    .D(net204),
    .Q(\clk_div.clock_sel_r ));
 sky130_fd_sc_hd__dfxtp_1 _2739_ (.CLK(clknet_4_2_0_net190),
    .D(_0049_),
    .Q(\wb_cross_clk.m_s_sync.d_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2740_ (.CLK(clknet_4_9_0_net190),
    .D(_0050_),
    .Q(\wb_cross_clk.m_s_sync.d_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2741_ (.CLK(clknet_4_2_0_net190),
    .D(_0051_),
    .Q(\wb_cross_clk.m_s_sync.d_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2742_ (.CLK(clknet_4_2_0_net190),
    .D(_0052_),
    .Q(\wb_cross_clk.m_s_sync.d_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2743_ (.CLK(clknet_4_3_0_net190),
    .D(_0053_),
    .Q(\wb_cross_clk.m_s_sync.d_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2744_ (.CLK(clknet_4_3_0_net190),
    .D(_0054_),
    .Q(\wb_cross_clk.m_s_sync.d_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2745_ (.CLK(clknet_4_0_0_net190),
    .D(_0055_),
    .Q(\wb_cross_clk.m_s_sync.d_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2746_ (.CLK(clknet_4_0_0_net190),
    .D(_0056_),
    .Q(\wb_cross_clk.m_s_sync.d_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2747_ (.CLK(clknet_4_3_0_net190),
    .D(_0057_),
    .Q(\wb_cross_clk.m_s_sync.d_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2748_ (.CLK(clknet_4_3_0_net190),
    .D(_0058_),
    .Q(\wb_cross_clk.m_s_sync.d_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2749_ (.CLK(clknet_4_6_0_net190),
    .D(_0059_),
    .Q(\wb_cross_clk.m_s_sync.d_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2750_ (.CLK(clknet_4_13_0_net190),
    .D(_0060_),
    .Q(\wb_cross_clk.m_s_sync.d_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2751_ (.CLK(clknet_4_6_0_net190),
    .D(_0061_),
    .Q(\wb_cross_clk.m_s_sync.d_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2752_ (.CLK(clknet_4_3_0_net190),
    .D(_0062_),
    .Q(\wb_cross_clk.m_s_sync.d_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2753_ (.CLK(clknet_4_6_0_net190),
    .D(_0063_),
    .Q(\wb_cross_clk.m_s_sync.d_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2754_ (.CLK(clknet_4_7_0_net190),
    .D(_0064_),
    .Q(\wb_cross_clk.m_s_sync.d_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2755_ (.CLK(clknet_4_6_0_net190),
    .D(_0065_),
    .Q(\wb_cross_clk.m_s_sync.d_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2756_ (.CLK(clknet_4_6_0_net190),
    .D(_0066_),
    .Q(\wb_cross_clk.m_s_sync.d_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2757_ (.CLK(clknet_4_7_0_net190),
    .D(_0067_),
    .Q(\wb_cross_clk.m_s_sync.d_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2758_ (.CLK(clknet_4_6_0_net190),
    .D(_0068_),
    .Q(\wb_cross_clk.m_s_sync.d_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2759_ (.CLK(clknet_4_7_0_net190),
    .D(_0069_),
    .Q(\wb_cross_clk.m_s_sync.d_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2760_ (.CLK(clknet_4_6_0_net190),
    .D(_0070_),
    .Q(\wb_cross_clk.m_s_sync.d_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2761_ (.CLK(clknet_4_1_0_net190),
    .D(_0071_),
    .Q(\wb_cross_clk.m_s_sync.d_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2762_ (.CLK(clknet_4_7_0_net190),
    .D(_0072_),
    .Q(\wb_cross_clk.m_s_sync.d_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2763_ (.CLK(clknet_4_1_0_net190),
    .D(_0073_),
    .Q(\wb_cross_clk.m_s_sync.d_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2764_ (.CLK(clknet_4_1_0_net190),
    .D(_0074_),
    .Q(\wb_cross_clk.m_s_sync.d_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2765_ (.CLK(clknet_4_4_0_net190),
    .D(_0075_),
    .Q(\wb_cross_clk.m_s_sync.d_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2766_ (.CLK(clknet_4_4_0_net190),
    .D(_0076_),
    .Q(\wb_cross_clk.m_s_sync.d_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2767_ (.CLK(clknet_4_4_0_net190),
    .D(_0077_),
    .Q(\wb_cross_clk.m_s_sync.d_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2768_ (.CLK(clknet_4_4_0_net190),
    .D(_0078_),
    .Q(\wb_cross_clk.m_s_sync.d_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2769_ (.CLK(clknet_4_4_0_net190),
    .D(_0079_),
    .Q(\wb_cross_clk.m_s_sync.d_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2770_ (.CLK(clknet_4_4_0_net190),
    .D(_0080_),
    .Q(\wb_cross_clk.m_s_sync.d_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2771_ (.CLK(clknet_4_4_0_net190),
    .D(_0081_),
    .Q(\wb_cross_clk.m_s_sync.d_data[32] ));
 sky130_fd_sc_hd__dfxtp_1 _2772_ (.CLK(clknet_4_4_0_net190),
    .D(_0082_),
    .Q(\wb_cross_clk.m_s_sync.d_data[33] ));
 sky130_fd_sc_hd__dfxtp_1 _2773_ (.CLK(clknet_4_5_0_net190),
    .D(_0083_),
    .Q(\wb_cross_clk.m_s_sync.d_data[34] ));
 sky130_fd_sc_hd__dfxtp_1 _2774_ (.CLK(clknet_4_5_0_net190),
    .D(_0084_),
    .Q(\wb_cross_clk.m_s_sync.d_data[35] ));
 sky130_fd_sc_hd__dfxtp_1 _2775_ (.CLK(clknet_4_5_0_net190),
    .D(_0085_),
    .Q(\wb_cross_clk.m_s_sync.d_data[36] ));
 sky130_fd_sc_hd__dfxtp_1 _2776_ (.CLK(clknet_4_4_0_net190),
    .D(_0086_),
    .Q(\wb_cross_clk.m_s_sync.d_data[37] ));
 sky130_fd_sc_hd__dfxtp_1 _2777_ (.CLK(clknet_4_5_0_net190),
    .D(_0087_),
    .Q(\wb_cross_clk.m_s_sync.d_data[38] ));
 sky130_fd_sc_hd__dfxtp_1 _2778_ (.CLK(clknet_4_5_0_net190),
    .D(_0088_),
    .Q(\wb_cross_clk.m_s_sync.d_data[39] ));
 sky130_fd_sc_hd__dfxtp_1 _2779_ (.CLK(clknet_4_5_0_net190),
    .D(_0089_),
    .Q(\wb_cross_clk.m_s_sync.d_data[40] ));
 sky130_fd_sc_hd__dfxtp_1 _2780_ (.CLK(clknet_4_5_0_net190),
    .D(_0090_),
    .Q(\wb_cross_clk.m_s_sync.d_data[41] ));
 sky130_fd_sc_hd__dfxtp_1 _2781_ (.CLK(clknet_4_5_0_net190),
    .D(_0091_),
    .Q(\wb_cross_clk.m_s_sync.d_data[42] ));
 sky130_fd_sc_hd__dfxtp_1 _2782_ (.CLK(clknet_4_5_0_net190),
    .D(_0092_),
    .Q(\wb_cross_clk.m_s_sync.d_data[43] ));
 sky130_fd_sc_hd__dfxtp_1 _2783_ (.CLK(clknet_4_7_0_net190),
    .D(_0093_),
    .Q(\wb_cross_clk.m_s_sync.d_data[44] ));
 sky130_fd_sc_hd__dfxtp_1 _2784_ (.CLK(clknet_4_5_0_net190),
    .D(_0094_),
    .Q(\wb_cross_clk.m_s_sync.d_data[45] ));
 sky130_fd_sc_hd__dfxtp_1 _2785_ (.CLK(clknet_4_0_0_net190),
    .D(_0095_),
    .Q(\wb_cross_clk.m_s_sync.d_data[46] ));
 sky130_fd_sc_hd__dfxtp_1 _2786_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0096_),
    .Q(\wb_cross_clk.prev_ack ));
 sky130_fd_sc_hd__dfxtp_1 _2787_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0097_),
    .Q(\wb_cross_clk.m_s_sync.s_xfer_xor_flag ));
 sky130_fd_sc_hd__dfxtp_1 _2788_ (.CLK(clknet_4_0_0_net190),
    .D(net425),
    .Q(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2789_ (.CLK(clknet_4_0_0_net190),
    .D(_0099_),
    .Q(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2790_ (.CLK(clknet_4_0_0_net190),
    .D(_0100_),
    .Q(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2791_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0101_),
    .Q(\wb_cross_clk.msy_xor_ack ));
 sky130_fd_sc_hd__dfxtp_1 _2792_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0102_),
    .Q(\wb_cross_clk.msy_xor_err ));
 sky130_fd_sc_hd__dfxtp_1 _2793_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0103_),
    .Q(\wb_cross_clk.m_wb_i_dat[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2794_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0104_),
    .Q(\wb_cross_clk.m_wb_i_dat[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2795_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0105_),
    .Q(\wb_cross_clk.m_wb_i_dat[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2796_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0106_),
    .Q(\wb_cross_clk.m_wb_i_dat[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2797_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0107_),
    .Q(\wb_cross_clk.m_wb_i_dat[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2798_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0108_),
    .Q(\wb_cross_clk.m_wb_i_dat[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2799_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0109_),
    .Q(\wb_cross_clk.m_wb_i_dat[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2800_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0110_),
    .Q(\wb_cross_clk.m_wb_i_dat[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2801_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0111_),
    .Q(\wb_cross_clk.m_wb_i_dat[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2802_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0112_),
    .Q(\wb_cross_clk.m_wb_i_dat[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2803_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0113_),
    .Q(\wb_cross_clk.m_wb_i_dat[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2804_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0114_),
    .Q(\wb_cross_clk.m_wb_i_dat[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2805_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0115_),
    .Q(\wb_cross_clk.m_wb_i_dat[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2806_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0116_),
    .Q(\wb_cross_clk.m_wb_i_dat[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2807_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0117_),
    .Q(\wb_cross_clk.m_wb_i_dat[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2808_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0118_),
    .Q(\wb_cross_clk.m_wb_i_dat[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2809_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0119_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2810_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0120_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2811_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0121_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2812_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0122_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2813_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0123_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2814_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0124_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2815_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0125_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2816_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0126_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2817_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0127_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2818_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0128_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2819_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0129_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2820_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0130_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2821_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0131_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2822_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0132_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2823_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0133_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2824_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0134_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2825_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0135_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2826_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0136_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2827_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0137_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2828_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0138_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2829_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0139_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2830_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0140_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2831_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0141_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2832_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0142_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2833_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0143_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2834_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0144_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2835_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0145_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2836_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0146_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2837_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0147_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2838_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0148_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2839_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0149_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2840_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0150_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2841_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0151_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[32] ));
 sky130_fd_sc_hd__dfxtp_1 _2842_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0152_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[33] ));
 sky130_fd_sc_hd__dfxtp_1 _2843_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0153_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[34] ));
 sky130_fd_sc_hd__dfxtp_1 _2844_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0154_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[35] ));
 sky130_fd_sc_hd__dfxtp_1 _2845_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0155_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[36] ));
 sky130_fd_sc_hd__dfxtp_1 _2846_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0156_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[37] ));
 sky130_fd_sc_hd__dfxtp_1 _2847_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0157_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[38] ));
 sky130_fd_sc_hd__dfxtp_1 _2848_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0158_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[39] ));
 sky130_fd_sc_hd__dfxtp_1 _2849_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0159_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[40] ));
 sky130_fd_sc_hd__dfxtp_1 _2850_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0160_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[41] ));
 sky130_fd_sc_hd__dfxtp_1 _2851_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0161_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[42] ));
 sky130_fd_sc_hd__dfxtp_1 _2852_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0162_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[43] ));
 sky130_fd_sc_hd__dfxtp_1 _2853_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0163_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[44] ));
 sky130_fd_sc_hd__dfxtp_1 _2854_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0164_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[45] ));
 sky130_fd_sc_hd__dfxtp_1 _2855_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0165_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[46] ));
 sky130_fd_sc_hd__dfxtp_1 _2856_ (.CLK(clknet_4_3_0_net190),
    .D(_0166_),
    .Q(\wb_cross_clk.s_m_sync.s_xfer_xor_flag ));
 sky130_fd_sc_hd__dfxtp_1 _2857_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0167_),
    .Q(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2858_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0168_),
    .Q(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2859_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0169_),
    .Q(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2860_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0170_),
    .Q(\wb_cross_clk.prev_stb ));
 sky130_fd_sc_hd__dfxtp_1 _2861_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0171_),
    .Q(\wb_cross_clk.prev_xor_err ));
 sky130_fd_sc_hd__dfxtp_1 _2862_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0172_),
    .Q(\wb_cross_clk.m_new_req_flag ));
 sky130_fd_sc_hd__dfxtp_1 _2863_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0173_),
    .Q(\wb_cross_clk.m_burst_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2864_ (.CLK(clknet_leaf_3_user_clock2),
    .D(net710),
    .Q(\wb_cross_clk.m_burst_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2865_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0175_),
    .Q(\wb_cross_clk.m_burst_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2866_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0176_),
    .Q(\wb_cross_clk.m_burst_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2867_ (.CLK(clknet_4_9_0_net190),
    .D(net567),
    .Q(\wb_cross_clk.s_burst_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2868_ (.CLK(clknet_4_9_0_net190),
    .D(net574),
    .Q(\wb_cross_clk.s_burst_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2869_ (.CLK(clknet_4_9_0_net190),
    .D(net593),
    .Q(\wb_cross_clk.s_burst_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2870_ (.CLK(clknet_4_9_0_net190),
    .D(_0180_),
    .Q(\wb_cross_clk.s_burst_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2871_ (.CLK(clknet_4_9_0_net190),
    .D(_0181_),
    .Q(\wb_cross_clk.ack_next_hold ));
 sky130_fd_sc_hd__dfxtp_1 _2872_ (.CLK(clknet_4_2_0_net190),
    .D(_0182_),
    .Q(\wb_cross_clk.err_xor_flag ));
 sky130_fd_sc_hd__dfxtp_1 _2873_ (.CLK(clknet_4_2_0_net190),
    .D(_0183_),
    .Q(\wb_cross_clk.ack_xor_flag ));
 sky130_fd_sc_hd__dfxtp_1 _2874_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0184_),
    .Q(\wb_cross_clk.prev_xor_ack ));
 sky130_fd_sc_hd__dfxtp_1 _2875_ (.CLK(clknet_4_9_0_net190),
    .D(_0185_),
    .Q(\wb_cross_clk.prev_xor_newreq ));
 sky130_fd_sc_hd__dfxtp_1 _2876_ (.CLK(clknet_4_12_0_net190),
    .D(_0186_),
    .Q(\wb_compressor.l_we ));
 sky130_fd_sc_hd__dfxtp_1 _2877_ (.CLK(clknet_4_12_0_net190),
    .D(_0187_),
    .Q(\wb_compressor.burst_end[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2878_ (.CLK(clknet_4_13_0_net190),
    .D(_0188_),
    .Q(\wb_compressor.burst_end[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2879_ (.CLK(clknet_4_12_0_net190),
    .D(_0189_),
    .Q(\wb_compressor.burst_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2880_ (.CLK(clknet_4_13_0_net190),
    .D(_0190_),
    .Q(\wb_compressor.burst_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2881_ (.CLK(clknet_4_14_0_net190),
    .D(net722),
    .Q(\wb_compressor.burst_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2882_ (.CLK(clknet_4_10_0_net190),
    .D(_0192_),
    .Q(\wb_compressor.wb_i_dat[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2883_ (.CLK(clknet_4_10_0_net190),
    .D(_0193_),
    .Q(\wb_compressor.wb_i_dat[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2884_ (.CLK(clknet_4_10_0_net190),
    .D(_0194_),
    .Q(\wb_compressor.wb_i_dat[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2885_ (.CLK(clknet_4_10_0_net190),
    .D(_0195_),
    .Q(\wb_compressor.wb_i_dat[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2886_ (.CLK(clknet_4_10_0_net190),
    .D(_0196_),
    .Q(\wb_compressor.wb_i_dat[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2887_ (.CLK(clknet_4_10_0_net190),
    .D(_0197_),
    .Q(\wb_compressor.wb_i_dat[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2888_ (.CLK(clknet_4_10_0_net190),
    .D(_0198_),
    .Q(\wb_compressor.wb_i_dat[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2889_ (.CLK(clknet_4_11_0_net190),
    .D(_0199_),
    .Q(\wb_compressor.wb_i_dat[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2890_ (.CLK(clknet_4_14_0_net190),
    .D(_0200_),
    .Q(\wb_compressor.wb_i_dat[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2891_ (.CLK(clknet_4_15_0_net190),
    .D(_0201_),
    .Q(\wb_compressor.wb_i_dat[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2892_ (.CLK(clknet_4_15_0_net190),
    .D(_0202_),
    .Q(\wb_compressor.wb_i_dat[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2893_ (.CLK(clknet_4_15_0_net190),
    .D(_0203_),
    .Q(\wb_compressor.wb_i_dat[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2894_ (.CLK(clknet_4_15_0_net190),
    .D(_0204_),
    .Q(\wb_compressor.wb_i_dat[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2895_ (.CLK(clknet_4_15_0_net190),
    .D(_0205_),
    .Q(\wb_compressor.wb_i_dat[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2896_ (.CLK(clknet_4_15_0_net190),
    .D(_0206_),
    .Q(\wb_compressor.wb_i_dat[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2897_ (.CLK(clknet_4_14_0_net190),
    .D(_0207_),
    .Q(\wb_compressor.wb_i_dat[15] ));
 sky130_fd_sc_hd__dfxtp_2 _2898_ (.CLK(clknet_4_11_0_net190),
    .D(net918),
    .Q(\wb_compressor.wb_ack ));
 sky130_fd_sc_hd__dfxtp_1 _2899_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0209_),
    .Q(\sspi.sy_clk[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2900_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0210_),
    .Q(\sspi.sy_clk[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2901_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0211_),
    .Q(\sspi.sy_clk[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2902_ (.CLK(clknet_4_11_0_net190),
    .D(net646),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_1 _2903_ (.CLK(clknet_4_11_0_net190),
    .D(_0213_),
    .Q(net199));
 sky130_fd_sc_hd__dfxtp_1 _2904_ (.CLK(clknet_4_8_0_net190),
    .D(net662),
    .Q(net173));
 sky130_fd_sc_hd__dfxtp_1 _2905_ (.CLK(clknet_4_8_0_net190),
    .D(net629),
    .Q(net174));
 sky130_fd_sc_hd__dfxtp_1 _2906_ (.CLK(clknet_4_8_0_net190),
    .D(net619),
    .Q(net175));
 sky130_fd_sc_hd__dfxtp_1 _2907_ (.CLK(clknet_4_8_0_net190),
    .D(net599),
    .Q(net176));
 sky130_fd_sc_hd__dfxtp_1 _2908_ (.CLK(clknet_4_8_0_net190),
    .D(net656),
    .Q(net177));
 sky130_fd_sc_hd__dfxtp_1 _2909_ (.CLK(clknet_4_8_0_net190),
    .D(net683),
    .Q(net178));
 sky130_fd_sc_hd__dfxtp_1 _2910_ (.CLK(clknet_4_8_0_net190),
    .D(net651),
    .Q(net179));
 sky130_fd_sc_hd__dfxtp_1 _2911_ (.CLK(clknet_4_8_0_net190),
    .D(net643),
    .Q(net180));
 sky130_fd_sc_hd__dfxtp_1 _2912_ (.CLK(clknet_4_8_0_net190),
    .D(net609),
    .Q(net181));
 sky130_fd_sc_hd__dfxtp_1 _2913_ (.CLK(clknet_4_8_0_net190),
    .D(net624),
    .Q(net182));
 sky130_fd_sc_hd__dfxtp_1 _2914_ (.CLK(clknet_4_8_0_net190),
    .D(net586),
    .Q(net184));
 sky130_fd_sc_hd__dfxtp_1 _2915_ (.CLK(clknet_4_8_0_net190),
    .D(net591),
    .Q(net185));
 sky130_fd_sc_hd__dfxtp_1 _2916_ (.CLK(clknet_4_9_0_net190),
    .D(net614),
    .Q(net186));
 sky130_fd_sc_hd__dfxtp_1 _2917_ (.CLK(clknet_4_9_0_net190),
    .D(net571),
    .Q(net187));
 sky130_fd_sc_hd__dfxtp_1 _2918_ (.CLK(clknet_4_9_0_net190),
    .D(net604),
    .Q(net188));
 sky130_fd_sc_hd__dfxtp_1 _2919_ (.CLK(clknet_4_9_0_net190),
    .D(net581),
    .Q(net189));
 sky130_fd_sc_hd__dfxtp_1 _2920_ (.CLK(clknet_4_12_0_net190),
    .D(net639),
    .Q(\wb_compressor.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2921_ (.CLK(clknet_4_14_0_net190),
    .D(_0000_),
    .Q(\wb_compressor.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2922_ (.CLK(clknet_4_12_0_net190),
    .D(_0011_),
    .Q(\wb_compressor.state[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2923_ (.CLK(clknet_4_12_0_net190),
    .D(_0001_),
    .Q(\wb_compressor.state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2924_ (.CLK(clknet_4_14_0_net190),
    .D(net670),
    .Q(\wb_compressor.state[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2925_ (.CLK(clknet_4_14_0_net190),
    .D(net691),
    .Q(\wb_compressor.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2926_ (.CLK(clknet_4_12_0_net190),
    .D(_0014_),
    .Q(\wb_compressor.state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2927_ (.CLK(clknet_leaf_28_user_clock2),
    .D(net870),
    .Q(\sspi.state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2928_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0003_),
    .Q(\sspi.state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2929_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0004_),
    .Q(\sspi.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2930_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0005_),
    .Q(\sspi.state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2931_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0006_),
    .Q(\sspi.state[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2932_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0007_),
    .Q(\sspi.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2933_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0008_),
    .Q(\sspi.state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2934_ (.CLK(clknet_leaf_4_user_clock2),
    .D(net699),
    .Q(\sspi.state[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2935_ (.CLK(clknet_leaf_32_user_clock2),
    .D(net689),
    .Q(\sspi.resp_err ));
 sky130_fd_sc_hd__dfxtp_1 _2936_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0231_),
    .Q(\sspi.bit_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2937_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0232_),
    .Q(\sspi.bit_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2938_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0233_),
    .Q(\sspi.bit_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2939_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0234_),
    .Q(\sspi.bit_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2940_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0235_),
    .Q(\sspi.bit_cnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2941_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0236_),
    .Q(\sspi.res_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2942_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0237_),
    .Q(\sspi.res_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2943_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0238_),
    .Q(\sspi.res_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2944_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0239_),
    .Q(\sspi.res_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2945_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0240_),
    .Q(\sspi.res_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2946_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0241_),
    .Q(\sspi.res_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2947_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0242_),
    .Q(\sspi.res_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2948_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0243_),
    .Q(\sspi.res_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2949_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0244_),
    .Q(\sspi.res_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2950_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0245_),
    .Q(\sspi.res_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2951_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0246_),
    .Q(\sspi.res_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2952_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0247_),
    .Q(\sspi.res_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2953_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0248_),
    .Q(\sspi.res_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2954_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0249_),
    .Q(\sspi.res_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2955_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0250_),
    .Q(\sspi.res_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2956_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0251_),
    .Q(\sspi.res_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2957_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0252_),
    .Q(\sspi.req_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2958_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0253_),
    .Q(\sspi.req_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2959_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0254_),
    .Q(\sspi.req_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2960_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0255_),
    .Q(\sspi.req_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2961_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0256_),
    .Q(\sspi.req_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2962_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0257_),
    .Q(\sspi.req_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2963_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0258_),
    .Q(\sspi.req_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2964_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0259_),
    .Q(\sspi.req_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2965_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0260_),
    .Q(\sspi.req_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2966_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0261_),
    .Q(\sspi.req_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2967_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0262_),
    .Q(\sspi.req_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2968_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0263_),
    .Q(\sspi.req_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2969_ (.CLK(clknet_leaf_25_user_clock2),
    .D(net701),
    .Q(\sspi.req_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2970_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0265_),
    .Q(\sspi.req_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2971_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0266_),
    .Q(\sspi.req_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2972_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0267_),
    .Q(\sspi.req_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2973_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0268_),
    .Q(\sspi.req_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2974_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0269_),
    .Q(\sspi.req_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2975_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0270_),
    .Q(\sspi.req_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2976_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0271_),
    .Q(\sspi.req_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2977_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0272_),
    .Q(\sspi.req_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2978_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0273_),
    .Q(\sspi.req_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2979_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0274_),
    .Q(\sspi.req_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2980_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0275_),
    .Q(\sspi.req_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2981_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0276_),
    .Q(\sspi.req_addr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2982_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0277_),
    .Q(\sspi.req_addr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2983_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0278_),
    .Q(\sspi.req_addr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2984_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0279_),
    .Q(\sspi.req_addr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2985_ (.CLK(clknet_leaf_25_user_clock2),
    .D(net693),
    .Q(\sspi.req_addr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2986_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0281_),
    .Q(\sspi.req_addr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2987_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0282_),
    .Q(\sspi.req_addr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2988_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0283_),
    .Q(\sspi.req_addr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2989_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0284_),
    .Q(\sspi.req_addr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2990_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0285_),
    .Q(\sspi.req_addr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2991_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0286_),
    .Q(\sspi.req_addr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2992_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0287_),
    .Q(\sspi.req_addr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2993_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0288_),
    .Q(\sspi.req_addr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2994_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0289_),
    .Q(\sspi.req_addr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2995_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0290_),
    .Q(\sspi.req_addr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2996_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0291_),
    .Q(\sspi.req_addr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2997_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0292_),
    .Q(\m_arbiter.wb0_adr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2998_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0293_),
    .Q(\m_arbiter.wb0_adr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2999_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0294_),
    .Q(\m_arbiter.wb0_adr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3000_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0295_),
    .Q(\m_arbiter.wb0_adr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3001_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0296_),
    .Q(\m_arbiter.wb0_adr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3002_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0297_),
    .Q(\m_arbiter.wb0_adr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3003_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0298_),
    .Q(\m_arbiter.wb0_adr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3004_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0299_),
    .Q(\m_arbiter.wb0_adr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3005_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0300_),
    .Q(\m_arbiter.wb0_adr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3006_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0301_),
    .Q(\m_arbiter.wb0_adr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3007_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0302_),
    .Q(\m_arbiter.wb0_adr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3008_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0303_),
    .Q(\m_arbiter.wb0_adr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3009_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0304_),
    .Q(\m_arbiter.wb0_adr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3010_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0305_),
    .Q(\m_arbiter.wb0_adr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3011_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0306_),
    .Q(\m_arbiter.wb0_adr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3012_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0307_),
    .Q(\m_arbiter.wb0_adr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3013_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0308_),
    .Q(\m_arbiter.wb0_adr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3014_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0309_),
    .Q(\m_arbiter.wb0_adr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3015_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0310_),
    .Q(\m_arbiter.wb0_adr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3016_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0311_),
    .Q(\m_arbiter.wb0_adr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3017_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0312_),
    .Q(\m_arbiter.wb0_adr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3018_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0313_),
    .Q(\m_arbiter.wb0_adr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3019_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0314_),
    .Q(\m_arbiter.wb0_adr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3020_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0315_),
    .Q(\m_arbiter.wb0_adr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3021_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0316_),
    .Q(\m_arbiter.wb0_we ));
 sky130_fd_sc_hd__dfxtp_1 _3022_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0317_),
    .Q(\m_arbiter.wb0_o_dat[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3023_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0318_),
    .Q(\m_arbiter.wb0_o_dat[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3024_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0319_),
    .Q(\m_arbiter.wb0_o_dat[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3025_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0320_),
    .Q(\m_arbiter.wb0_o_dat[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3026_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0321_),
    .Q(\m_arbiter.wb0_o_dat[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3027_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0322_),
    .Q(\m_arbiter.wb0_o_dat[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3028_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0323_),
    .Q(\m_arbiter.wb0_o_dat[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3029_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0324_),
    .Q(\m_arbiter.wb0_o_dat[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3030_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0325_),
    .Q(\m_arbiter.wb0_o_dat[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3031_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0326_),
    .Q(\m_arbiter.wb0_o_dat[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3032_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0327_),
    .Q(\m_arbiter.wb0_o_dat[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3033_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0328_),
    .Q(\m_arbiter.wb0_o_dat[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3034_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0329_),
    .Q(\m_arbiter.wb0_o_dat[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3035_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0330_),
    .Q(\m_arbiter.wb0_o_dat[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3036_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0331_),
    .Q(\m_arbiter.wb0_o_dat[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3037_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0332_),
    .Q(\m_arbiter.wb0_o_dat[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3038_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0333_),
    .Q(\clk_div.cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3039_ (.CLK(clknet_leaf_36_user_clock2),
    .D(net882),
    .Q(\clk_div.cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3040_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0335_),
    .Q(\clk_div.cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3041_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0336_),
    .Q(\clk_div.cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3042_ (.CLK(clknet_leaf_36_user_clock2),
    .D(net697),
    .Q(\clk_div.cnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3043_ (.CLK(clknet_leaf_36_user_clock2),
    .D(_0338_),
    .Q(\clk_div.cnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3044_ (.CLK(clknet_leaf_36_user_clock2),
    .D(_0339_),
    .Q(\clk_div.cnt[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3045_ (.CLK(clknet_leaf_36_user_clock2),
    .D(net736),
    .Q(\clk_div.cnt[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3046_ (.CLK(clknet_leaf_36_user_clock2),
    .D(_0341_),
    .Q(\clk_div.cnt[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3047_ (.CLK(clknet_leaf_1_user_clock2),
    .D(net731),
    .Q(\clk_div.cnt[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3048_ (.CLK(clknet_leaf_1_user_clock2),
    .D(net719),
    .Q(\clk_div.cnt[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3049_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0344_),
    .Q(\clk_div.cnt[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3050_ (.CLK(clknet_leaf_1_user_clock2),
    .D(net713),
    .Q(\clk_div.cnt[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3051_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0346_),
    .Q(\clk_div.cnt[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3052_ (.CLK(clknet_leaf_1_user_clock2),
    .D(net727),
    .Q(\clk_div.cnt[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3053_ (.CLK(clknet_leaf_1_user_clock2),
    .D(net695),
    .Q(\clk_div.cnt[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3054_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0349_),
    .Q(\m_arbiter.i_wb0_cyc ));
 sky130_fd_sc_hd__dfxtp_2 _3055_ (.CLK(clknet_leaf_4_user_clock2),
    .D(net864),
    .Q(net193));
 sky130_fd_sc_hd__dfxtp_2 _3056_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0351_),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_2 _3057_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0352_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_2 _3058_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0353_),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_2 _3059_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0354_),
    .Q(net167));
 sky130_fd_sc_hd__dfxtp_2 _3060_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0355_),
    .Q(net168));
 sky130_fd_sc_hd__dfxtp_2 _3061_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0356_),
    .Q(net169));
 sky130_fd_sc_hd__dfxtp_2 _3062_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0357_),
    .Q(net170));
 sky130_fd_sc_hd__dfxtp_2 _3063_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0358_),
    .Q(net171));
 sky130_fd_sc_hd__dfxtp_2 _3064_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0359_),
    .Q(net172));
 sky130_fd_sc_hd__dfxtp_2 _3065_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0360_),
    .Q(net183));
 sky130_fd_sc_hd__dfxtp_2 _3066_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0361_),
    .Q(net192));
 sky130_fd_sc_hd__dfxtp_2 _3067_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0362_),
    .Q(net194));
 sky130_fd_sc_hd__dfxtp_2 _3068_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0363_),
    .Q(net195));
 sky130_fd_sc_hd__dfxtp_2 _3069_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0364_),
    .Q(net196));
 sky130_fd_sc_hd__dfxtp_2 _3070_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0365_),
    .Q(net197));
 sky130_fd_sc_hd__dfxtp_2 _3071_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0366_),
    .Q(net198));
 sky130_fd_sc_hd__dfstp_1 _3072_ (.CLK(clknet_leaf_10_user_clock2),
    .D(net206),
    .SET_B(_0015_),
    .Q(\rst_soc_sync.reset_sync_ff[0] ));
 sky130_fd_sc_hd__dfstp_4 _3073_ (.CLK(clknet_leaf_11_user_clock2),
    .D(net672),
    .SET_B(_0016_),
    .Q(net103));
 sky130_fd_sc_hd__dfstp_1 _3074_ (.CLK(clknet_4_10_0_net190),
    .D(net205),
    .SET_B(net754),
    .Q(\rst_cw_sync.reset_sync_ff[0] ));
 sky130_fd_sc_hd__dfstp_1 _3075_ (.CLK(clknet_4_11_0_net190),
    .D(net671),
    .SET_B(net831),
    .Q(net191));
 sky130_fd_sc_hd__dfxtp_1 _3076_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0367_),
    .Q(\m_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__conb_1 interconnect_outer_414 (.HI(net414));
 sky130_fd_sc_hd__conb_1 interconnect_outer_415 (.HI(net415));
 sky130_fd_sc_hd__conb_1 interconnect_outer_416 (.HI(net416));
 sky130_fd_sc_hd__conb_1 interconnect_outer_417 (.HI(net417));
 sky130_fd_sc_hd__conb_1 interconnect_outer_418 (.HI(net418));
 sky130_fd_sc_hd__conb_1 interconnect_outer_419 (.HI(net419));
 sky130_fd_sc_hd__conb_1 interconnect_outer_420 (.HI(net420));
 sky130_fd_sc_hd__conb_1 interconnect_outer_421 (.HI(net421));
 sky130_fd_sc_hd__conb_1 interconnect_outer_422 (.HI(net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_0_user_clock2));
 sky130_fd_sc_hd__conb_1 _3072__206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 interconnect_outer_207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 interconnect_outer_208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 interconnect_outer_209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 interconnect_outer_210 (.LO(net210));
 sky130_fd_sc_hd__conb_1 interconnect_outer_211 (.LO(net211));
 sky130_fd_sc_hd__conb_1 interconnect_outer_212 (.LO(net212));
 sky130_fd_sc_hd__conb_1 interconnect_outer_213 (.LO(net213));
 sky130_fd_sc_hd__conb_1 interconnect_outer_214 (.LO(net214));
 sky130_fd_sc_hd__conb_1 interconnect_outer_215 (.LO(net215));
 sky130_fd_sc_hd__conb_1 interconnect_outer_216 (.LO(net216));
 sky130_fd_sc_hd__conb_1 interconnect_outer_217 (.LO(net217));
 sky130_fd_sc_hd__conb_1 interconnect_outer_218 (.LO(net218));
 sky130_fd_sc_hd__conb_1 interconnect_outer_219 (.LO(net219));
 sky130_fd_sc_hd__conb_1 interconnect_outer_220 (.LO(net220));
 sky130_fd_sc_hd__conb_1 interconnect_outer_221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 interconnect_outer_222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 interconnect_outer_223 (.LO(net223));
 sky130_fd_sc_hd__conb_1 interconnect_outer_224 (.LO(net224));
 sky130_fd_sc_hd__conb_1 interconnect_outer_225 (.LO(net225));
 sky130_fd_sc_hd__conb_1 interconnect_outer_226 (.LO(net226));
 sky130_fd_sc_hd__conb_1 interconnect_outer_227 (.LO(net227));
 sky130_fd_sc_hd__conb_1 interconnect_outer_228 (.LO(net228));
 sky130_fd_sc_hd__conb_1 interconnect_outer_229 (.LO(net229));
 sky130_fd_sc_hd__conb_1 interconnect_outer_230 (.LO(net230));
 sky130_fd_sc_hd__conb_1 interconnect_outer_231 (.LO(net231));
 sky130_fd_sc_hd__conb_1 interconnect_outer_232 (.LO(net232));
 sky130_fd_sc_hd__conb_1 interconnect_outer_233 (.LO(net233));
 sky130_fd_sc_hd__conb_1 interconnect_outer_234 (.LO(net234));
 sky130_fd_sc_hd__conb_1 interconnect_outer_235 (.LO(net235));
 sky130_fd_sc_hd__conb_1 interconnect_outer_236 (.LO(net236));
 sky130_fd_sc_hd__conb_1 interconnect_outer_237 (.LO(net237));
 sky130_fd_sc_hd__conb_1 interconnect_outer_238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 interconnect_outer_239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 interconnect_outer_240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 interconnect_outer_241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 interconnect_outer_242 (.LO(net242));
 sky130_fd_sc_hd__conb_1 interconnect_outer_243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 interconnect_outer_244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 interconnect_outer_245 (.LO(net245));
 sky130_fd_sc_hd__conb_1 interconnect_outer_246 (.LO(net246));
 sky130_fd_sc_hd__conb_1 interconnect_outer_247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 interconnect_outer_248 (.LO(net248));
 sky130_fd_sc_hd__conb_1 interconnect_outer_249 (.LO(net249));
 sky130_fd_sc_hd__conb_1 interconnect_outer_250 (.LO(net250));
 sky130_fd_sc_hd__conb_1 interconnect_outer_251 (.LO(net251));
 sky130_fd_sc_hd__conb_1 interconnect_outer_252 (.LO(net252));
 sky130_fd_sc_hd__conb_1 interconnect_outer_253 (.LO(net253));
 sky130_fd_sc_hd__conb_1 interconnect_outer_254 (.LO(net254));
 sky130_fd_sc_hd__conb_1 interconnect_outer_255 (.LO(net255));
 sky130_fd_sc_hd__conb_1 interconnect_outer_256 (.LO(net256));
 sky130_fd_sc_hd__conb_1 interconnect_outer_257 (.LO(net257));
 sky130_fd_sc_hd__conb_1 interconnect_outer_258 (.LO(net258));
 sky130_fd_sc_hd__conb_1 interconnect_outer_259 (.LO(net259));
 sky130_fd_sc_hd__conb_1 interconnect_outer_260 (.LO(net260));
 sky130_fd_sc_hd__conb_1 interconnect_outer_261 (.LO(net261));
 sky130_fd_sc_hd__conb_1 interconnect_outer_262 (.LO(net262));
 sky130_fd_sc_hd__conb_1 interconnect_outer_263 (.LO(net263));
 sky130_fd_sc_hd__conb_1 interconnect_outer_264 (.LO(net264));
 sky130_fd_sc_hd__conb_1 interconnect_outer_265 (.LO(net265));
 sky130_fd_sc_hd__conb_1 interconnect_outer_266 (.LO(net266));
 sky130_fd_sc_hd__conb_1 interconnect_outer_267 (.LO(net267));
 sky130_fd_sc_hd__conb_1 interconnect_outer_268 (.LO(net268));
 sky130_fd_sc_hd__conb_1 interconnect_outer_269 (.LO(net269));
 sky130_fd_sc_hd__conb_1 interconnect_outer_270 (.LO(net270));
 sky130_fd_sc_hd__conb_1 interconnect_outer_271 (.LO(net271));
 sky130_fd_sc_hd__conb_1 interconnect_outer_272 (.LO(net272));
 sky130_fd_sc_hd__conb_1 interconnect_outer_273 (.LO(net273));
 sky130_fd_sc_hd__conb_1 interconnect_outer_274 (.LO(net274));
 sky130_fd_sc_hd__conb_1 interconnect_outer_275 (.LO(net275));
 sky130_fd_sc_hd__conb_1 interconnect_outer_276 (.LO(net276));
 sky130_fd_sc_hd__conb_1 interconnect_outer_277 (.LO(net277));
 sky130_fd_sc_hd__conb_1 interconnect_outer_278 (.LO(net278));
 sky130_fd_sc_hd__conb_1 interconnect_outer_279 (.LO(net279));
 sky130_fd_sc_hd__conb_1 interconnect_outer_280 (.LO(net280));
 sky130_fd_sc_hd__conb_1 interconnect_outer_281 (.LO(net281));
 sky130_fd_sc_hd__conb_1 interconnect_outer_282 (.LO(net282));
 sky130_fd_sc_hd__conb_1 interconnect_outer_283 (.LO(net283));
 sky130_fd_sc_hd__conb_1 interconnect_outer_284 (.LO(net284));
 sky130_fd_sc_hd__conb_1 interconnect_outer_285 (.LO(net285));
 sky130_fd_sc_hd__conb_1 interconnect_outer_286 (.LO(net286));
 sky130_fd_sc_hd__conb_1 interconnect_outer_287 (.LO(net287));
 sky130_fd_sc_hd__conb_1 interconnect_outer_288 (.LO(net288));
 sky130_fd_sc_hd__conb_1 interconnect_outer_289 (.LO(net289));
 sky130_fd_sc_hd__conb_1 interconnect_outer_290 (.LO(net290));
 sky130_fd_sc_hd__conb_1 interconnect_outer_291 (.LO(net291));
 sky130_fd_sc_hd__conb_1 interconnect_outer_292 (.LO(net292));
 sky130_fd_sc_hd__conb_1 interconnect_outer_293 (.LO(net293));
 sky130_fd_sc_hd__conb_1 interconnect_outer_294 (.LO(net294));
 sky130_fd_sc_hd__conb_1 interconnect_outer_295 (.LO(net295));
 sky130_fd_sc_hd__conb_1 interconnect_outer_296 (.LO(net296));
 sky130_fd_sc_hd__conb_1 interconnect_outer_297 (.LO(net297));
 sky130_fd_sc_hd__conb_1 interconnect_outer_298 (.LO(net298));
 sky130_fd_sc_hd__conb_1 interconnect_outer_299 (.LO(net299));
 sky130_fd_sc_hd__conb_1 interconnect_outer_300 (.LO(net300));
 sky130_fd_sc_hd__conb_1 interconnect_outer_301 (.LO(net301));
 sky130_fd_sc_hd__conb_1 interconnect_outer_302 (.LO(net302));
 sky130_fd_sc_hd__conb_1 interconnect_outer_303 (.LO(net303));
 sky130_fd_sc_hd__conb_1 interconnect_outer_304 (.LO(net304));
 sky130_fd_sc_hd__conb_1 interconnect_outer_305 (.LO(net305));
 sky130_fd_sc_hd__conb_1 interconnect_outer_306 (.LO(net306));
 sky130_fd_sc_hd__conb_1 interconnect_outer_307 (.LO(net307));
 sky130_fd_sc_hd__conb_1 interconnect_outer_308 (.LO(net308));
 sky130_fd_sc_hd__conb_1 interconnect_outer_309 (.LO(net309));
 sky130_fd_sc_hd__conb_1 interconnect_outer_310 (.LO(net310));
 sky130_fd_sc_hd__conb_1 interconnect_outer_311 (.LO(net311));
 sky130_fd_sc_hd__conb_1 interconnect_outer_312 (.LO(net312));
 sky130_fd_sc_hd__conb_1 interconnect_outer_313 (.LO(net313));
 sky130_fd_sc_hd__conb_1 interconnect_outer_314 (.LO(net314));
 sky130_fd_sc_hd__conb_1 interconnect_outer_315 (.LO(net315));
 sky130_fd_sc_hd__conb_1 interconnect_outer_316 (.LO(net316));
 sky130_fd_sc_hd__conb_1 interconnect_outer_317 (.LO(net317));
 sky130_fd_sc_hd__conb_1 interconnect_outer_318 (.LO(net318));
 sky130_fd_sc_hd__conb_1 interconnect_outer_319 (.LO(net319));
 sky130_fd_sc_hd__conb_1 interconnect_outer_320 (.LO(net320));
 sky130_fd_sc_hd__conb_1 interconnect_outer_321 (.LO(net321));
 sky130_fd_sc_hd__conb_1 interconnect_outer_322 (.LO(net322));
 sky130_fd_sc_hd__conb_1 interconnect_outer_323 (.LO(net323));
 sky130_fd_sc_hd__conb_1 interconnect_outer_324 (.LO(net324));
 sky130_fd_sc_hd__conb_1 interconnect_outer_325 (.LO(net325));
 sky130_fd_sc_hd__conb_1 interconnect_outer_326 (.LO(net326));
 sky130_fd_sc_hd__conb_1 interconnect_outer_327 (.LO(net327));
 sky130_fd_sc_hd__conb_1 interconnect_outer_328 (.LO(net328));
 sky130_fd_sc_hd__conb_1 interconnect_outer_329 (.LO(net329));
 sky130_fd_sc_hd__conb_1 interconnect_outer_330 (.LO(net330));
 sky130_fd_sc_hd__conb_1 interconnect_outer_331 (.LO(net331));
 sky130_fd_sc_hd__conb_1 interconnect_outer_332 (.LO(net332));
 sky130_fd_sc_hd__conb_1 interconnect_outer_333 (.LO(net333));
 sky130_fd_sc_hd__conb_1 interconnect_outer_334 (.LO(net334));
 sky130_fd_sc_hd__conb_1 interconnect_outer_335 (.LO(net335));
 sky130_fd_sc_hd__conb_1 interconnect_outer_336 (.LO(net336));
 sky130_fd_sc_hd__conb_1 interconnect_outer_337 (.LO(net337));
 sky130_fd_sc_hd__conb_1 interconnect_outer_338 (.LO(net338));
 sky130_fd_sc_hd__conb_1 interconnect_outer_339 (.LO(net339));
 sky130_fd_sc_hd__conb_1 interconnect_outer_340 (.LO(net340));
 sky130_fd_sc_hd__conb_1 interconnect_outer_341 (.LO(net341));
 sky130_fd_sc_hd__conb_1 interconnect_outer_342 (.LO(net342));
 sky130_fd_sc_hd__conb_1 interconnect_outer_343 (.LO(net343));
 sky130_fd_sc_hd__conb_1 interconnect_outer_344 (.LO(net344));
 sky130_fd_sc_hd__conb_1 interconnect_outer_345 (.LO(net345));
 sky130_fd_sc_hd__conb_1 interconnect_outer_346 (.LO(net346));
 sky130_fd_sc_hd__conb_1 interconnect_outer_347 (.LO(net347));
 sky130_fd_sc_hd__conb_1 interconnect_outer_348 (.LO(net348));
 sky130_fd_sc_hd__conb_1 interconnect_outer_349 (.LO(net349));
 sky130_fd_sc_hd__conb_1 interconnect_outer_350 (.LO(net350));
 sky130_fd_sc_hd__conb_1 interconnect_outer_351 (.LO(net351));
 sky130_fd_sc_hd__conb_1 interconnect_outer_352 (.LO(net352));
 sky130_fd_sc_hd__conb_1 interconnect_outer_353 (.LO(net353));
 sky130_fd_sc_hd__conb_1 interconnect_outer_354 (.LO(net354));
 sky130_fd_sc_hd__conb_1 interconnect_outer_355 (.LO(net355));
 sky130_fd_sc_hd__conb_1 interconnect_outer_356 (.LO(net356));
 sky130_fd_sc_hd__conb_1 interconnect_outer_357 (.LO(net357));
 sky130_fd_sc_hd__conb_1 interconnect_outer_358 (.LO(net358));
 sky130_fd_sc_hd__conb_1 interconnect_outer_359 (.LO(net359));
 sky130_fd_sc_hd__conb_1 interconnect_outer_360 (.LO(net360));
 sky130_fd_sc_hd__conb_1 interconnect_outer_361 (.LO(net361));
 sky130_fd_sc_hd__conb_1 interconnect_outer_362 (.LO(net362));
 sky130_fd_sc_hd__conb_1 interconnect_outer_363 (.LO(net363));
 sky130_fd_sc_hd__conb_1 interconnect_outer_364 (.LO(net364));
 sky130_fd_sc_hd__conb_1 interconnect_outer_365 (.LO(net365));
 sky130_fd_sc_hd__conb_1 interconnect_outer_366 (.LO(net366));
 sky130_fd_sc_hd__conb_1 interconnect_outer_367 (.LO(net367));
 sky130_fd_sc_hd__conb_1 interconnect_outer_368 (.LO(net368));
 sky130_fd_sc_hd__conb_1 interconnect_outer_369 (.LO(net369));
 sky130_fd_sc_hd__conb_1 interconnect_outer_370 (.LO(net370));
 sky130_fd_sc_hd__conb_1 interconnect_outer_371 (.LO(net371));
 sky130_fd_sc_hd__conb_1 interconnect_outer_372 (.LO(net372));
 sky130_fd_sc_hd__conb_1 interconnect_outer_373 (.LO(net373));
 sky130_fd_sc_hd__conb_1 interconnect_outer_374 (.LO(net374));
 sky130_fd_sc_hd__conb_1 interconnect_outer_375 (.LO(net375));
 sky130_fd_sc_hd__conb_1 interconnect_outer_376 (.LO(net376));
 sky130_fd_sc_hd__conb_1 interconnect_outer_377 (.LO(net377));
 sky130_fd_sc_hd__conb_1 interconnect_outer_378 (.LO(net378));
 sky130_fd_sc_hd__conb_1 interconnect_outer_379 (.LO(net379));
 sky130_fd_sc_hd__conb_1 interconnect_outer_380 (.LO(net380));
 sky130_fd_sc_hd__conb_1 interconnect_outer_381 (.LO(net381));
 sky130_fd_sc_hd__conb_1 interconnect_outer_382 (.LO(net382));
 sky130_fd_sc_hd__conb_1 interconnect_outer_383 (.LO(net383));
 sky130_fd_sc_hd__conb_1 interconnect_outer_384 (.LO(net384));
 sky130_fd_sc_hd__conb_1 interconnect_outer_385 (.LO(net385));
 sky130_fd_sc_hd__conb_1 interconnect_outer_386 (.LO(net386));
 sky130_fd_sc_hd__conb_1 interconnect_outer_387 (.LO(net387));
 sky130_fd_sc_hd__conb_1 interconnect_outer_388 (.LO(net388));
 sky130_fd_sc_hd__conb_1 interconnect_outer_389 (.LO(net389));
 sky130_fd_sc_hd__conb_1 interconnect_outer_390 (.LO(net390));
 sky130_fd_sc_hd__conb_1 interconnect_outer_391 (.LO(net391));
 sky130_fd_sc_hd__conb_1 interconnect_outer_392 (.LO(net392));
 sky130_fd_sc_hd__conb_1 interconnect_outer_393 (.LO(net393));
 sky130_fd_sc_hd__conb_1 interconnect_outer_394 (.LO(net394));
 sky130_fd_sc_hd__conb_1 interconnect_outer_395 (.LO(net395));
 sky130_fd_sc_hd__conb_1 interconnect_outer_396 (.LO(net396));
 sky130_fd_sc_hd__conb_1 interconnect_outer_397 (.LO(net397));
 sky130_fd_sc_hd__conb_1 interconnect_outer_398 (.LO(net398));
 sky130_fd_sc_hd__conb_1 interconnect_outer_399 (.LO(net399));
 sky130_fd_sc_hd__conb_1 interconnect_outer_400 (.LO(net400));
 sky130_fd_sc_hd__conb_1 interconnect_outer_401 (.LO(net401));
 sky130_fd_sc_hd__conb_1 interconnect_outer_402 (.LO(net402));
 sky130_fd_sc_hd__conb_1 interconnect_outer_403 (.LO(net403));
 sky130_fd_sc_hd__conb_1 interconnect_outer_404 (.LO(net404));
 sky130_fd_sc_hd__conb_1 interconnect_outer_405 (.LO(net405));
 sky130_fd_sc_hd__conb_1 interconnect_outer_406 (.LO(net406));
 sky130_fd_sc_hd__conb_1 interconnect_outer_407 (.LO(net407));
 sky130_fd_sc_hd__conb_1 interconnect_outer_408 (.LO(net408));
 sky130_fd_sc_hd__conb_1 interconnect_outer_409 (.LO(net409));
 sky130_fd_sc_hd__conb_1 interconnect_outer_410 (.LO(net410));
 sky130_fd_sc_hd__conb_1 interconnect_outer_411 (.LO(net411));
 sky130_fd_sc_hd__conb_1 interconnect_outer_412 (.LO(net412));
 sky130_fd_sc_hd__conb_1 interconnect_outer_413 (.HI(net413));
 sky130_fd_sc_hd__buf_2 _3295_ (.A(clknet_opt_1_0_user_clock2),
    .X(net99));
 sky130_fd_sc_hd__buf_2 _3296_ (.A(clknet_opt_2_0_user_clock2),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 _3297_ (.A(net202),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _3298_ (.A(net202),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 _3299_ (.A(net202),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 _3300_ (.A(net202),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 _3301_ (.A(net202),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 _3302_ (.A(net202),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 _3303_ (.A(net202),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 _3304_ (.A(net202),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 _3305_ (.A(net202),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 _3306_ (.A(net203),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 _3307_ (.A(net203),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 _3308_ (.A(net203),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 _3309_ (.A(net203),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 _3310_ (.A(net203),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 _3311_ (.A(net203),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 _3312_ (.A(net202),
    .X(net200));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(inner_wb_4_burst),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(inner_wb_8_burst),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(inner_wb_adr[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(inner_wb_adr[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(inner_wb_adr[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(inner_wb_adr[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(inner_wb_adr[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(inner_wb_adr[14]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(inner_wb_adr[15]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(inner_wb_adr[16]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(inner_wb_adr[17]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(inner_wb_adr[18]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(inner_wb_adr[19]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(inner_wb_adr[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(inner_wb_adr[20]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(inner_wb_adr[21]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(inner_wb_adr[22]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(inner_wb_adr[23]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(inner_wb_adr[2]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(inner_wb_adr[3]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(inner_wb_adr[4]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(inner_wb_adr[5]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(inner_wb_adr[6]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(inner_wb_adr[7]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(inner_wb_adr[8]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(inner_wb_adr[9]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(inner_wb_cyc),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(inner_wb_o_dat[0]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(inner_wb_o_dat[10]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(inner_wb_o_dat[11]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(inner_wb_o_dat[12]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(inner_wb_o_dat[13]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(inner_wb_o_dat[14]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(inner_wb_o_dat[15]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(inner_wb_o_dat[1]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(inner_wb_o_dat[2]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(inner_wb_o_dat[3]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(inner_wb_o_dat[4]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(inner_wb_o_dat[5]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(inner_wb_o_dat[6]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(inner_wb_o_dat[7]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(inner_wb_o_dat[8]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(inner_wb_o_dat[9]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(inner_wb_sel[0]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(inner_wb_sel[1]),
    .X(net45));
 sky130_fd_sc_hd__dlymetal6s2s_1 input46 (.A(inner_wb_stb),
    .X(net46));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(inner_wb_we),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(iram_o_data[0]),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(iram_o_data[10]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(iram_o_data[11]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(iram_o_data[12]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(iram_o_data[13]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(iram_o_data[14]),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 input54 (.A(iram_o_data[15]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(iram_o_data[1]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(iram_o_data[2]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(iram_o_data[3]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(iram_o_data[4]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(iram_o_data[5]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(iram_o_data[6]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(iram_o_data[7]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(iram_o_data[8]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(iram_o_data[9]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(net753),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(la_oenb[0]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(m_io_in[0]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(m_io_in[10]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(m_io_in[11]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(m_io_in[12]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(m_io_in[13]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(m_io_in[14]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(m_io_in[15]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(m_io_in[16]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(m_io_in[17]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(m_io_in[18]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(m_io_in[19]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(m_io_in[1]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(m_io_in[20]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(m_io_in[21]),
    .X(net79));
 sky130_fd_sc_hd__dlymetal6s2s_1 input80 (.A(m_io_in[22]),
    .X(net80));
 sky130_fd_sc_hd__dlymetal6s2s_1 input81 (.A(m_io_in[23]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(m_io_in[24]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(m_io_in[25]),
    .X(net83));
 sky130_fd_sc_hd__buf_2 input84 (.A(m_io_in[26]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(m_io_in[27]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(m_io_in[2]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(m_io_in[30]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(m_io_in[31]),
    .X(net88));
 sky130_fd_sc_hd__buf_2 input89 (.A(m_io_in[32]),
    .X(net89));
 sky130_fd_sc_hd__buf_4 input90 (.A(m_io_in[33]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 input91 (.A(m_io_in[34]),
    .X(net91));
 sky130_fd_sc_hd__buf_4 input92 (.A(m_io_in[35]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(m_io_in[3]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(m_io_in[4]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(m_io_in[5]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(m_io_in[6]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(m_io_in[7]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(net830),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net99),
    .X(inner_clock));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(inner_disable));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(inner_embed_mode));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(inner_ext_irq));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(inner_reset));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(inner_wb_ack));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(inner_wb_err));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(inner_wb_i_dat[0]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(inner_wb_i_dat[10]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(inner_wb_i_dat[11]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(inner_wb_i_dat[12]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(inner_wb_i_dat[13]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(inner_wb_i_dat[14]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(inner_wb_i_dat[15]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(inner_wb_i_dat[1]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(inner_wb_i_dat[2]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(inner_wb_i_dat[3]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(inner_wb_i_dat[4]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(inner_wb_i_dat[5]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(inner_wb_i_dat[6]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(inner_wb_i_dat[7]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(inner_wb_i_dat[8]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(inner_wb_i_dat[9]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(iram_addr[0]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(iram_addr[1]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(iram_addr[2]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(iram_addr[3]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(iram_addr[4]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(iram_addr[5]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(iram_addr[6]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(iram_addr[7]));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net130),
    .X(iram_clk));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(iram_i_data[0]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(iram_i_data[10]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(iram_i_data[11]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(iram_i_data[12]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(iram_i_data[13]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(iram_i_data[14]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(iram_i_data[15]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(iram_i_data[1]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(iram_i_data[2]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(iram_i_data[3]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(iram_i_data[4]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(iram_i_data[5]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(iram_i_data[6]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(iram_i_data[7]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(iram_i_data[8]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(iram_i_data[9]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(iram_we));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(m_io_oeb[0]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(m_io_oeb[10]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(m_io_oeb[11]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(m_io_oeb[12]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(m_io_oeb[13]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(m_io_oeb[14]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(m_io_oeb[15]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(m_io_oeb[16]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(m_io_oeb[17]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(m_io_oeb[18]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(m_io_oeb[19]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(m_io_oeb[1]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(m_io_oeb[20]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(m_io_oeb[21]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(m_io_oeb[22]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(m_io_oeb[23]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(m_io_oeb[24]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net203),
    .X(m_io_oeb[25]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(m_io_oeb[2]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(m_io_oeb[3]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(m_io_oeb[4]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(m_io_oeb[5]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(m_io_oeb[6]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(m_io_oeb[7]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(m_io_out[0]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(m_io_out[10]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(m_io_out[11]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(m_io_out[12]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(m_io_out[13]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(m_io_out[14]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(m_io_out[15]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(m_io_out[16]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(m_io_out[17]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(m_io_out[18]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(m_io_out[19]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(m_io_out[1]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(m_io_out[20]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(m_io_out[21]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(m_io_out[22]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(m_io_out[23]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(m_io_out[24]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(m_io_out[25]));
 sky130_fd_sc_hd__clkbuf_1 output190 (.A(clknet_4_10_0_net190),
    .X(m_io_out[28]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(m_io_out[29]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(m_io_out[2]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(m_io_out[36]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(m_io_out[3]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(m_io_out[4]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(m_io_out[5]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(m_io_out[6]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(m_io_out[7]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(m_io_out[8]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(m_io_out[9]));
 sky130_fd_sc_hd__clkbuf_4 fanout201 (.A(net191),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 fanout203 (.A(net165),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(net568),
    .X(net204));
 sky130_fd_sc_hd__conb_1 _3074__205 (.LO(net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_1_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_2_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_3_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_5_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_6_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_7_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_8_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_10_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_12_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_13_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_14_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_16_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_17_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_20_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_22_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_23_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_24_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_25_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_26_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_27_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_28_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_29_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_30_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_33_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_34_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_36_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_user_clock2 (.A(user_clock2),
    .X(clknet_0_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_opt_1_0_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_opt_2_0_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net190 (.A(net190),
    .X(clknet_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_0_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_1_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_2_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_3_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_4_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_5_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_6_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_7_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_8_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_9_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_10_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_11_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_12_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_13_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_14_0_net190));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_net190 (.A(clknet_0_net190),
    .X(clknet_4_15_0_net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\wb_cross_clk.m_s_sync.s_xfer_xor_flag ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0661_),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0098_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\wb_cross_clk.m_s_sync.s_data_ff[27] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0610_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0611_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\wb_cross_clk.m_s_sync.s_data_ff[12] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0578_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0579_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\wb_cross_clk.m_s_sync.s_data_ff[10] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0574_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0575_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\wb_cross_clk.m_s_sync.s_data_ff[17] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0588_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0589_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\wb_cross_clk.m_s_sync.s_data_ff[14] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0582_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0583_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\wb_cross_clk.m_s_sync.s_data_ff[1] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0554_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0555_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\wb_cross_clk.m_s_sync.s_data_ff[26] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0608_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0609_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\wb_cross_clk.m_s_sync.s_data_ff[8] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0569_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0570_),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\wb_cross_clk.m_s_sync.s_data_ff[16] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_0586_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0587_),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\wb_cross_clk.m_s_sync.s_data_ff[5] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0562_),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_0563_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\wb_cross_clk.m_s_sync.s_data_ff[45] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_0649_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0650_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\wb_cross_clk.m_s_sync.s_data_ff[43] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0645_),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0646_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\wb_cross_clk.m_s_sync.s_data_ff[11] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0576_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0577_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\wb_cross_clk.m_s_sync.s_data_ff[19] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0593_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0594_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\wb_cross_clk.m_s_sync.s_data_ff[13] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0580_),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0581_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\wb_cross_clk.m_s_sync.s_data_ff[7] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0566_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0567_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\wb_cross_clk.m_s_sync.s_data_ff[18] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0591_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0592_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\wb_cross_clk.m_s_sync.s_data_ff[25] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0606_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0607_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\wb_cross_clk.m_s_sync.s_data_ff[23] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0602_),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0603_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\wb_cross_clk.m_s_sync.s_data_ff[34] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0626_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0627_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\wb_cross_clk.m_s_sync.s_data_ff[21] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0598_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0599_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\wb_cross_clk.m_s_sync.s_data_ff[6] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0564_),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0565_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\wb_cross_clk.m_s_sync.s_data_ff[9] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0571_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0572_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\wb_cross_clk.m_s_sync.s_data_ff[20] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0596_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0597_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\wb_cross_clk.m_s_sync.s_data_ff[24] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0604_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0605_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\wb_cross_clk.m_s_sync.s_data_ff[33] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0624_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_0625_),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\wb_cross_clk.m_s_sync.s_data_ff[3] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_0558_),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0559_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\wb_cross_clk.m_s_sync.s_data_ff[15] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0584_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_0585_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\wb_cross_clk.m_s_sync.s_data_ff[37] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0632_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0633_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\wb_cross_clk.m_s_sync.s_data_ff[40] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0639_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0640_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\wb_cross_clk.m_s_sync.s_data_ff[0] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0552_),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0553_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\wb_cross_clk.m_s_sync.s_data_ff[44] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0647_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0648_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\wb_cross_clk.m_s_sync.s_data_ff[41] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0641_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0642_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\wb_cross_clk.m_s_sync.s_data_ff[4] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0560_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0561_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\wb_cross_clk.m_s_sync.s_data_ff[31] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0620_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0621_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\wb_cross_clk.m_s_sync.s_data_ff[29] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0615_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0616_),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\wb_cross_clk.m_s_sync.s_data_ff[2] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0556_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_0557_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\wb_cross_clk.m_s_sync.s_data_ff[22] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0600_),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0601_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\wb_cross_clk.m_s_sync.s_data_ff[42] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0643_),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0644_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\wb_cross_clk.m_s_sync.s_data_ff[32] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0622_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0623_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\wb_cross_clk.m_s_sync.s_data_ff[39] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_0637_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0638_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\wb_cross_clk.m_s_sync.s_data_ff[30] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0618_),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0619_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\wb_cross_clk.m_s_sync.s_data_ff[28] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_0613_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0614_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\wb_cross_clk.m_s_sync.s_data_ff[46] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0651_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0652_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\wb_cross_clk.m_s_sync.s_data_ff[38] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0635_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\wb_cross_clk.m_s_sync.s_data_ff[35] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0628_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\wb_cross_clk.m_s_sync.s_data_ff[36] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0630_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\m_arbiter.wb0_we ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0479_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0791_),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0177_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\clk_div.clock_sel ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_1325_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0923_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0227_),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\wb_cross_clk.s_burst_cnt[1] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0793_),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0178_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\wb_compressor.l_we ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0811_),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\m_arbiter.wb0_adr[15] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_1261_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_1319_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0929_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_0229_),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\m_arbiter.wb0_adr[18] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_1246_),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_1320_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_0912_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0224_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\m_arbiter.wb0_adr[19] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_1248_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_1323_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0916_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_0225_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\wb_cross_clk.s_burst_cnt[2] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_0179_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\m_arbiter.wb0_o_dat[3] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_1231_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0882_),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_0883_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0884_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0217_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\m_arbiter.wb0_adr[14] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_1260_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_1321_),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0926_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0228_),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\m_arbiter.wb0_adr[16] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_1249_),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_1324_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_0904_),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0222_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\m_arbiter.wb0_adr[20] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_1252_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_1318_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0920_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0226_),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\m_arbiter.wb0_o_dat[2] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_1232_),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_0876_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0880_),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_0216_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\m_arbiter.wb0_adr[17] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_1247_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_1314_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_0908_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0223_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\m_arbiter.wb0_adr[1] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_1238_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0868_),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_0874_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0215_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\m_arbiter.wb0_adr[22] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_1254_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0481_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_0482_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\m_arbiter.wb0_adr[21] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_1253_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_1276_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_1288_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_0369_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0010_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\m_arbiter.wb0_o_dat[7] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_0898_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_0900_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_0221_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(net165),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0849_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_0212_),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\m_arbiter.wb0_o_dat[6] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_1227_),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_0896_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0897_),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0220_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\m_arbiter.wb0_o_dat[4] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0886_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0887_),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0888_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_0218_),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\m_arbiter.wb0_adr[0] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_1240_),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0865_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0866_),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_0867_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0214_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\split_s_ff[0] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\disable_s_ff[0] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\irq_s_ff[0] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\wb_compressor.burst_end[2] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0816_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\wb_compressor.state[6] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_1306_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0012_),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\rst_cw_sync.reset_sync_ff[0] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\rst_soc_sync.reset_sync_ff[0] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\wb_compressor.wb_err ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_0019_),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\embed_s_ff[0] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\wb_compressor.burst_end[0] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0815_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\m_arbiter.wb0_o_dat[5] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_1228_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_0891_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_0892_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_0893_),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_0219_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(net199),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_0858_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\wb_cross_clk.s_m_sync.s_xfer_xor_flag ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\clk_div.res_clk ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\sspi.resp_err ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_0230_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\wb_compressor.state[2] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_0013_),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\sspi.req_addr[12] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_0280_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\clk_div.cnt[15] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0348_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\clk_div.cnt[4] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_0337_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\sspi.state[3] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_0009_),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\sspi.req_data[12] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_0264_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\sspi.state[6] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\clk_div.next_div_val ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0539_),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[0] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\sspi.req_data[9] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_1130_),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\wb_cross_clk.m_burst_cnt[0] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_0776_),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_0174_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\clk_div.cnt[12] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_1165_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_0345_),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\sspi.req_data[4] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\m_arbiter.i_wb0_cyc ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\sspi.req_addr[21] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\clk_div.cnt[10] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_1161_),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_0343_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\sspi.req_data[1] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\wb_compressor.burst_cnt[2] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_0191_),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[0] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\sspi.req_data[3] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\clk_div.cnt[14] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_1169_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(_0347_),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\sspi.sy_clk[0] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\clk_div.cnt[9] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_1159_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_0342_),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\clk_div.cnt[11] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\sspi.req_addr[9] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_1103_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\clk_div.cnt[7] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0340_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\m_arbiter.wb0_o_dat[8] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\clk_div.cnt[13] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\wb_cross_clk.s_m_sync.s_data_ff[12] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_0512_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\m_arbiter.wb0_adr[11] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\sspi.req_data[2] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\sspi.req_addr[4] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\wb_cross_clk.s_m_sync.s_data_ff[1] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_0500_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\sspi.req_data[15] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(_1136_),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\wb_cross_clk.s_m_sync.s_data_ff[7] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0507_),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\m_arbiter.wb0_adr[5] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\sspi.req_addr[7] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_1100_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(la_data_in[0]),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_0017_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\clk_div.cnt[6] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_1152_),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\wb_cross_clk.m_new_req_flag ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\sspi.req_addr[15] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\m_arbiter.wb0_o_dat[11] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\wb_cross_clk.s_m_sync.s_data_ff[14] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(_0514_),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\m_arbiter.wb0_o_dat[1] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\sspi.req_addr[13] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_1107_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\m_arbiter.wb0_adr[4] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\m_arbiter.wb0_o_dat[13] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\sspi.req_addr[8] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\wb_cross_clk.s_m_sync.s_data_ff[11] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(_0511_),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\sspi.req_data[7] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\m_arbiter.wb0_adr[23] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\sspi.req_addr[5] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\sspi.req_data[13] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_1134_),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\m_arbiter.wb0_o_dat[0] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\clk_div.next_div_buff[0] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\m_arbiter.wb0_o_dat[12] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\m_arbiter.wb0_o_dat[10] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(_1131_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\sspi.res_data[8] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\m_arbiter.wb0_adr[2] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(net103),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\sspi.bit_cnt[3] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\sspi.req_addr[0] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\sspi.req_data[14] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_1135_),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\m_arbiter.wb0_adr[12] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\sspi.req_addr[1] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\clk_div.next_div_buff[2] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\wb_cross_clk.s_m_sync.s_data_ff[8] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(_0508_),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\sspi.req_addr[19] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\sspi.req_addr[22] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\sspi.req_data[11] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(_1132_),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\sspi.state[1] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\sspi.req_data[5] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\sspi.req_addr[18] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\sspi.res_data[9] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\sspi.req_addr[14] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\wb_cross_clk.s_m_sync.s_data_ff[4] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_0503_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\sspi.bit_cnt[4] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_1045_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\sspi.req_addr[16] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\sspi.bit_cnt[2] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\sspi.bit_cnt[4] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\m_arbiter.wb0_adr[3] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(_1096_),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\sspi.res_data[4] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\m_arbiter.wb0_adr[8] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_1263_),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\sspi.req_data[6] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\wb_cross_clk.s_m_sync.s_data_ff[13] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(_0513_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\clk_div.next_div_buff[3] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\sspi.req_data[8] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\m_arbiter.wb0_adr[10] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\wb_cross_clk.s_m_sync.s_data_ff[5] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_0504_),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\sspi.bit_cnt[1] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_1006_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\sspi.res_data[5] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\sspi.req_addr[10] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\sspi.req_addr[23] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\sspi.state[4] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\sspi.req_data[10] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\wb_cross_clk.s_m_sync.s_data_ff[9] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(_0509_),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(mgt_wb_rst_i),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(_0018_),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\sspi.req_addr[2] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\sspi.req_addr[6] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_1099_),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\sspi.bit_cnt[2] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\m_arbiter.wb0_adr[13] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\sspi.res_data[6] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\wb_cross_clk.s_m_sync.s_data_ff[2] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(_0501_),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\wb_cross_clk.s_m_sync.s_data_ff[15] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(_0515_),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\sspi.state[2] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\clk_div.next_div_buff[1] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\sspi.res_data[7] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\wb_cross_clk.s_m_sync.s_data_ff[3] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0502_),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\wb_cross_clk.s_m_sync.s_data_ff[17] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0517_),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\sspi.req_addr[11] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\wb_cross_clk.s_m_sync.s_data_ff[16] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(_0516_),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\wb_cross_clk.s_m_sync.s_data_ff[10] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(_0510_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\sspi.req_addr[3] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\sspi.bit_cnt[0] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\wb_cross_clk.s_m_sync.s_data_ff[0] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(_0498_),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\wb_cross_clk.s_m_sync.s_data_ff[6] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(_0505_),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\sspi.res_data[10] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\sspi.req_addr[17] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\sspi.sy_clk[1] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(net193),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_0350_),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\sspi.state[7] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0402_),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\sspi.state[0] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\sspi.req_addr[20] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\sspi.state[5] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0002_),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\sspi.res_data[11] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\wb_cross_clk.m_s_sync.d_data[0] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\sspi.res_data[1] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\sspi.req_data[0] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\wb_cross_clk.s_burst_cnt[3] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\sspi.res_data[3] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\sspi.res_data[2] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\sspi.sy_clk[2] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\sspi.res_data[0] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\wb_compressor.wb_i_dat[11] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\clk_div.cnt[1] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_0334_),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\wb_cross_clk.ack_next_hold ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\wb_cross_clk.m_burst_cnt[3] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_0782_),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\sspi.res_data[12] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\wb_compressor.wb_i_dat[15] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\wb_compressor.wb_i_dat[7] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\sspi.res_data[13] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\wb_cross_clk.msy_xor_ack ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\wb_cross_clk.m_burst_cnt[2] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\wb_compressor.wb_i_dat[6] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\wb_cross_clk.msy_xor_err ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\wb_compressor.wb_i_dat[8] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\sspi.res_data[15] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\wb_compressor.wb_i_dat[2] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\wb_compressor.wb_i_dat[14] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\sspi.res_data[14] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\wb_compressor.wb_i_dat[5] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\wb_compressor.burst_cnt[1] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\wb_compressor.wb_i_dat[9] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\wb_compressor.wb_i_dat[13] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\wb_compressor.wb_i_dat[1] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(_0828_),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\wb_compressor.wb_i_dat[12] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\wb_cross_clk.prev_xor_ack ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_0653_),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\clk_div.curr_div[0] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\wb_compressor.wb_i_dat[10] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\wb_compressor.wb_i_dat[3] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_0830_),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\clk_div.curr_div[2] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\wb_compressor.wb_i_dat[0] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\wb_compressor.burst_cnt[0] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\wb_compressor.wb_ack ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_0208_),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\wb_cross_clk.m_wb_i_dat[8] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\wb_cross_clk.m_wb_i_dat[7] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\wb_cross_clk.m_wb_i_dat[13] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\wb_cross_clk.m_wb_i_dat[2] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\wb_cross_clk.m_wb_i_dat[12] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\wb_cross_clk.m_wb_i_dat[15] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\wb_cross_clk.m_wb_i_dat[5] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\wb_cross_clk.m_wb_i_dat[14] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\wb_cross_clk.m_wb_i_dat[4] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\wb_cross_clk.m_wb_i_dat[1] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\wb_cross_clk.m_wb_i_dat[10] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\wb_cross_clk.m_wb_i_dat[11] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\wb_cross_clk.m_wb_i_dat[3] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\clk_div.curr_div[3] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\wb_cross_clk.ack_xor_flag ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\wb_cross_clk.m_wb_i_dat[0] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\wb_cross_clk.m_wb_i_dat[6] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\wb_compressor.wb_i_dat[4] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\wb_cross_clk.m_wb_i_dat[9] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(net196),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\clk_div.cnt[5] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\clk_div.cnt[2] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(_1139_),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_1141_),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(net194),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\wb_cross_clk.err_xor_flag ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(_0499_),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\clk_div.cnt[3] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(_1144_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(net198),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\clk_div.cnt[0] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(net197),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(net172),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(net195),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(net192),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\clk_div.cnt[8] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(_1157_),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(net183),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\wb_compressor.state[4] ),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(net148),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(net169),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(net159),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(net171),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(net168),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(net167),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(net170),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(net166),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\sspi.state[1] ),
    .X(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold216_A (.DIODE(_0369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__A1 (.DIODE(_0369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2177__A1 (.DIODE(_0369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__A1 (.DIODE(_0369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__A (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__A (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__A (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__A (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2656__A (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__A (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__A (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__A (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1691__A (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__A (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__C (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2264__A1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__B (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1476__A1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2264__A2 (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1660__C (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__B (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1476__A2 (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2314__D (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__A (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2050__B1 (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2033__A (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__A (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__A (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1506__A (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1504__A (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1494__A (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__A1 (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2390__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1502__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__C1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__C1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__B (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__A (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__A (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__A (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2293__A1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__A (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__A (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__A2 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__A2 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__A2 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__A2 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__B (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__A (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__A (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__B (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__B (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__C (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__A (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2371__A (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__A (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__A (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2645__C1 (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__B1 (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__A1 (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2055__B1 (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__A (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__B1 (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__A (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__A (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__A (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__C1 (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__B1 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__C1 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__A (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1694__A (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__A1 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__A1 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1500__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1498__A (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__A1 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1515__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__A (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__A (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__A (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__A (.DIODE(_0423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1557__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1532__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__A (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2183__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1593__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__B1 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2040__B (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__B2 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1592__B2 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__B2 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__B2 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__B2 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__B2 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__B2 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__B2 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__B2 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2095__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__S (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__S (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1564__S (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1559__S (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1554__S (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1549__S (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__S (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__B1 (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__B1 (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1555__B1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__B1 (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1570__B1 (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__B1 (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1660__B (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1598__B (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__A2 (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1592__A2 (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__A2 (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__A2 (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__A2 (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__A2 (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__A2 (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__A2 (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__S (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__S (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2237__S (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__S (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2227__S (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__S (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__S (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__S (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__S (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__S (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__B1 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__B1 (.DIODE(_0471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__B1 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__B1 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__B1 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__B1 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1592__B1 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__B1 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold143_A (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__C (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2673__B (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__D (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__A1 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1678__C (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1598__C (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__A (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2137__S (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2135__S (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__S (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2131__S (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__S (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2127__S (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2125__S (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2123__S (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__B (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2083__A1 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2066__B1 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__B1 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1658__S (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__A (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__A (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__A2 (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2032__A2 (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2031__A2 (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__S (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__S (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__S (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__S (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__S (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__S (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__S (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1656__S (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1654__S (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__S (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1650__S (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1648__S (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__S (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__S (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__S (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__S (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__S (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__B1_N (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__B1_N (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__B (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__A2 (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1674__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__B (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1850__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1841__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1832__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__A (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__A (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__A (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1733__S (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1730__S (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1726__S (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__S (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1720__S (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__S (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1714__S (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1711__S (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1708__S (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__S (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1756__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1753__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1750__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1741__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1738__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1731__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1765__S (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1762__S (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__S (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1755__S (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__S (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1749__S (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__S (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__S (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__S (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1737__S (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1791__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1788__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1779__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1770__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1763__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1797__S (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__S (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1790__S (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__S (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__S (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__S (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__S (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__S (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__S (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__S (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1823__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1814__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1808__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1805__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1798__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1795__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1829__S (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1826__S (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1822__S (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__S (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1816__S (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__S (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__S (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__S (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1804__S (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1801__S (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__A (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1851__A (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__A (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1845__A (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1842__A (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__A (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__A (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1833__A (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1830__A (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1827__A (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2062__B1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__C1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2055__C1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__B (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__S (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__S (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__S (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__S (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__A2 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__A2 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1903__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1887__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2038__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1925__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1910__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1907__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1904__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2104__A0 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__A2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__C (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__A1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__A0 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__C (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__A0 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__A1 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2198__A0 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__A1 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2050__A1 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__B (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__B (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2025__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2004__A (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__A (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__A (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__A (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__S (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__S (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__S (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1954__S (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__S (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1950__S (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1948__S (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__S (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__S (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__S (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1996__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__S (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2021__S (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2019__S (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__S (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__S (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2013__S (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__S (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2009__S (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__S (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__S (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2300__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2159__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__B (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2042__B (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2040__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__B (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__S (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__S (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2223__S (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__S (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__S (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2208__S (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__S (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__S (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__S (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__S (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2261__A2 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__A2 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__A2 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__A3 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__A2 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2179__A (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2177__A2 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2173__C_N (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2249__B2 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__B2 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2239__B2 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__B2 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__A1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__A1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2243__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2198__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2221__A2 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2225__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__A2 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2239__A2 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__A2 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__S (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__S (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__S (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__S (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__S (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__S (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__A (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__D (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__A (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__A (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__S (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__S (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2499__S (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__S (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__S (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__S (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__S (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__S (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__A2 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__C1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__C1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2686__C1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__C1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__C1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__C1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__C1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__B1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__B1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__C1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__A2 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__B1 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__B1 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__B1 (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__D (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__B (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__B (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__C (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__A1 (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__A1 (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__A1 (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A1 (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__A (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__A (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2307__B (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__S (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2346__S (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__S (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__S (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__S (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__S (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__A (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2336__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A1 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2475__A2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__A2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__A1 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__A1 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__A0 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__A1 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__A0 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2368__A1 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__A0 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__B2 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__A2 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__A3 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A2 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2390__B (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__B (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__B (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__B (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold400_A (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__A2 (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__A2 (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__A2 (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__A2 (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__B (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2366__B (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__B (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__A (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__B (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__A (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__B (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A0 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__A0 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__A0 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__A0 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A0 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2426__A0 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2416__A0 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__A0 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__A0 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__A0 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold382_A (.DIODE(_1045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A0 (.DIODE(_1045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__A0 (.DIODE(_1045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__A0 (.DIODE(_1045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__A0 (.DIODE(_1045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__A0 (.DIODE(_1045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__A4 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__A2 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__A3 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__A4 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__A3 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__B (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__B (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__B (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__S (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__S (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__S (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__S (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__S (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__S (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__S (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__S (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__S (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__S (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__S (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__S (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__S (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__S (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2564__S (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__S (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__A (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__S (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__S (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__S (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__S (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__S (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__S (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2548__S (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__S (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__S (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__S (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1403__A1 (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1402__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1382__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1378__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1364__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1346__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1337__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1335__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1330__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__A1 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__A (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1933__A (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__A (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1514__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1512__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1510__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1342__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1333__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1332__A (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__A (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1597__S (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1524__S (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1522__S (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1520__S (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1518__S (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1516__S (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1344__S (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1340__S (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1338__S (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__S (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1373__S (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__S (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1368__S (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1367__S (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__S (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1360__S (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1353__S (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1351__S (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1349__S (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1387__S (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1386__S (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__S (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1384__S (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1381__S (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__S (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1375__S (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1370__S (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1369__S (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1356__S (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1361__A (.DIODE(_1242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1363__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold161_A (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__A1 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__A (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1371__A (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold199_A (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__A1 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__B (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1371__B (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__A1 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__A (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__A0 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1395__A_N (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1376__A (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold189_A (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2021__A1 (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__B (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1395__B (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1376__B (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold213_A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__B (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1376__C (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold209_A (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2025__A1 (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__D (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1376__D (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__A0 (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__A1 (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__C (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__A (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1379__A (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__A1 (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1450__A0 (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__C (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1383__A (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold179_A (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2009__A1 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1395__D (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1383__B (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold390_A (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2227__A0 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__A_N (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1388__A (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2237__A0 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__A1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__B (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1388__B (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__A0 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__A1 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__B (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1388__C (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__A0 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__A1 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__C (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1388__D (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold214_A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__B (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1473__B (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__B (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__A1 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1678__B (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1406__B (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__A2 (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1600__B1 (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1453__B1 (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__C (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1425__A2 (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__B1 (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1793__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1761__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1729__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1604__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1435__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2031__B1 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1721__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1718__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1712__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1709__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1706__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2262__A1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__A1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__A1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__A1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2225__B2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2221__A1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2209__A1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2204__A1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__A1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__A1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__A (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__A (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__A (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2081__A (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__A (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__A (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1436__A (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__C1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__C1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__C1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__C1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2201__C1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__C1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2186__C1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__C1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__B1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__B1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__S (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__S (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2104__S (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1543__A (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__A (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__S (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1446__S (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1441__S (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__S (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1439__S (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold200_A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__A (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold157_A (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__B (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold162_A (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__C (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold180_A (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__D (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold167_A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1452__A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold185_A (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1452__B (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold146_A (.DIODE(\clk_div.clock_sel ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(inner_wb_4_burst));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(inner_wb_8_burst));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(inner_wb_adr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(inner_wb_adr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(inner_wb_adr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(inner_wb_adr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(inner_wb_adr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(inner_wb_adr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(inner_wb_adr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(inner_wb_adr[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(inner_wb_adr[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(inner_wb_adr[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(inner_wb_adr[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(inner_wb_adr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(inner_wb_adr[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(inner_wb_adr[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(inner_wb_adr[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(inner_wb_adr[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(inner_wb_adr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(inner_wb_adr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(inner_wb_adr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(inner_wb_adr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(inner_wb_adr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(inner_wb_adr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(inner_wb_adr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(inner_wb_adr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(inner_wb_cyc));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(inner_wb_o_dat[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(inner_wb_o_dat[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(inner_wb_o_dat[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(inner_wb_o_dat[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(inner_wb_o_dat[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(inner_wb_o_dat[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(inner_wb_o_dat[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(inner_wb_o_dat[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(inner_wb_o_dat[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(inner_wb_o_dat[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(inner_wb_o_dat[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(inner_wb_o_dat[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(inner_wb_o_dat[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(inner_wb_o_dat[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(inner_wb_o_dat[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(inner_wb_o_dat[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(inner_wb_sel[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(inner_wb_sel[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(inner_wb_stb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(inner_wb_we));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(iram_o_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(iram_o_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(iram_o_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(iram_o_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(iram_o_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(iram_o_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(iram_o_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(iram_o_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(iram_o_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(iram_o_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(iram_o_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(iram_o_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(iram_o_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(iram_o_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(iram_o_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(iram_o_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold331_A (.DIODE(la_data_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(la_oenb[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(m_io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(m_io_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(m_io_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(m_io_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(m_io_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(m_io_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(m_io_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(m_io_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(m_io_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(m_io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(m_io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(m_io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(m_io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(m_io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(m_io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(m_io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(m_io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(m_io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(m_io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(m_io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(m_io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(m_io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(m_io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(m_io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(m_io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(m_io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(m_io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(m_io_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(m_io_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(m_io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(m_io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(m_io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold408_A (.DIODE(mgt_wb_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold413_A (.DIODE(\sspi.bit_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold384_A (.DIODE(\sspi.bit_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__B1 (.DIODE(\sspi.bit_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__C1 (.DIODE(\sspi.bit_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__A (.DIODE(\sspi.bit_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__A (.DIODE(\sspi.bit_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__A (.DIODE(\sspi.bit_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1480__A (.DIODE(\sspi.bit_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_user_clock2_A (.DIODE(user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2249__A1 (.DIODE(\wb_compressor.state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__A1 (.DIODE(\wb_compressor.state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2239__A1 (.DIODE(\wb_compressor.state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__A1 (.DIODE(\wb_compressor.state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__A1 (.DIODE(\wb_compressor.state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2199__A1 (.DIODE(\wb_compressor.state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__B2 (.DIODE(\wb_compressor.state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2097__A (.DIODE(\wb_compressor.state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1433__A (.DIODE(\wb_compressor.state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold495_A (.DIODE(\wb_compressor.wb_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__A (.DIODE(\wb_compressor.wb_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1472__A0 (.DIODE(\wb_compressor.wb_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1424__A (.DIODE(\wb_compressor.wb_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold251_A (.DIODE(\wb_compressor.wb_err ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__B (.DIODE(\wb_compressor.wb_err ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__B (.DIODE(\wb_compressor.wb_err ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__A0 (.DIODE(\wb_compressor.wb_err ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold514_A (.DIODE(\wb_compressor.wb_i_dat[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__A1 (.DIODE(\wb_compressor.wb_i_dat[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1559__A0 (.DIODE(\wb_compressor.wb_i_dat[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold462_A (.DIODE(\wb_cross_clk.ack_next_hold ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1407__A_N (.DIODE(\wb_cross_clk.ack_next_hold ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1356__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1378__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1382__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__1370__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__1367__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__1369__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__1373__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1375__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1518__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__1524__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1403__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__1597__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1592__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__1555__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__1570__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__1533__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2139__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2141__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2147__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2149__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2151__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__A_N (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1430__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1419__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__B2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__D (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__D (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__D (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__D_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1458__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__1490__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1558__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__2695__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__2694__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold360_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1492__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2346__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2336__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2183__A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1979__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1399__B_N (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1391__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1981__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__C_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1399__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1391__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__A0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1366__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1366__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__A0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1677__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1526__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1400__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__D_N (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__A0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__C (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__C (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1679__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__A0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__1967__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2243__A0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__A0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__1948__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1950__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1683__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2686__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2208__A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1954__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2223__A0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__A0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold536_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__1532__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold538_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold543_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold541_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1553__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold540_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__1557__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold537_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold542_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold539_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold529_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__1532__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_output173_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2186__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__2201__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_output176_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_output178_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_output180_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_output181_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2231__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_output182_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold534_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_output183_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_output184_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2241__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_output185_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_output186_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2251__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_output187_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_output188_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_output189_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2263__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net190_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold531_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_output192_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold441_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold521_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold530_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_output195_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__1557__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold516_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_output196_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold528_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_output197_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold526_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_output198_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold262_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_output199_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__1449__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__1448__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__1445__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__1444__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__1443__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__1472__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__D (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__1408__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__1438__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_1_0_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_2_0_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_net190_A (.DIODE(clknet_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__CLK (.DIODE(clknet_4_4_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__CLK (.DIODE(clknet_4_4_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__CLK (.DIODE(clknet_4_4_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__CLK (.DIODE(clknet_4_4_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__CLK (.DIODE(clknet_4_4_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__CLK (.DIODE(clknet_4_4_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__CLK (.DIODE(clknet_4_4_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__CLK (.DIODE(clknet_4_4_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__CLK (.DIODE(clknet_4_4_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__CLK (.DIODE(clknet_4_11_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2716__CLK (.DIODE(clknet_4_11_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__CLK (.DIODE(clknet_4_11_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__CLK (.DIODE(clknet_4_11_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2889__CLK (.DIODE(clknet_4_11_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2898__CLK (.DIODE(clknet_4_11_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2902__CLK (.DIODE(clknet_4_11_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2903__CLK (.DIODE(clknet_4_11_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__CLK (.DIODE(clknet_4_11_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2721__CLK (.DIODE(clknet_4_13_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2723__CLK (.DIODE(clknet_4_13_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__CLK (.DIODE(clknet_4_13_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2878__CLK (.DIODE(clknet_4_13_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__CLK (.DIODE(clknet_4_13_0_net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__A0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__2072__A (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__A (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1450__S (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__A (.DIODE(net917));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_622 ();
 assign iram1_addr[0] = net207;
 assign iram1_addr[1] = net208;
 assign iram1_addr[2] = net209;
 assign iram1_addr[3] = net210;
 assign iram1_addr[4] = net211;
 assign iram1_addr[5] = net212;
 assign iram1_addr[6] = net213;
 assign iram1_addr[7] = net214;
 assign iram_csb = net413;
 assign iram_i_data[16] = net215;
 assign iram_i_data[17] = net216;
 assign iram_i_data[18] = net217;
 assign iram_i_data[19] = net218;
 assign iram_i_data[20] = net219;
 assign iram_i_data[21] = net220;
 assign iram_i_data[22] = net221;
 assign iram_i_data[23] = net222;
 assign iram_i_data[24] = net223;
 assign iram_i_data[25] = net224;
 assign iram_i_data[26] = net225;
 assign iram_i_data[27] = net226;
 assign iram_i_data[28] = net227;
 assign iram_i_data[29] = net228;
 assign iram_i_data[30] = net229;
 assign iram_i_data[31] = net230;
 assign iram_w_mask[0] = net231;
 assign iram_w_mask[1] = net232;
 assign iram_w_mask[2] = net233;
 assign iram_w_mask[3] = net234;
 assign irq[0] = net235;
 assign irq[1] = net236;
 assign irq[2] = net237;
 assign la_data_out[0] = net238;
 assign la_data_out[100] = net338;
 assign la_data_out[101] = net339;
 assign la_data_out[102] = net340;
 assign la_data_out[103] = net341;
 assign la_data_out[104] = net342;
 assign la_data_out[105] = net343;
 assign la_data_out[106] = net344;
 assign la_data_out[107] = net345;
 assign la_data_out[108] = net346;
 assign la_data_out[109] = net347;
 assign la_data_out[10] = net248;
 assign la_data_out[110] = net348;
 assign la_data_out[111] = net349;
 assign la_data_out[112] = net350;
 assign la_data_out[113] = net351;
 assign la_data_out[114] = net352;
 assign la_data_out[115] = net353;
 assign la_data_out[116] = net354;
 assign la_data_out[117] = net355;
 assign la_data_out[118] = net356;
 assign la_data_out[119] = net357;
 assign la_data_out[11] = net249;
 assign la_data_out[120] = net358;
 assign la_data_out[121] = net359;
 assign la_data_out[122] = net360;
 assign la_data_out[123] = net361;
 assign la_data_out[124] = net362;
 assign la_data_out[125] = net363;
 assign la_data_out[126] = net364;
 assign la_data_out[127] = net365;
 assign la_data_out[12] = net250;
 assign la_data_out[13] = net251;
 assign la_data_out[14] = net252;
 assign la_data_out[15] = net253;
 assign la_data_out[16] = net254;
 assign la_data_out[17] = net255;
 assign la_data_out[18] = net256;
 assign la_data_out[19] = net257;
 assign la_data_out[1] = net239;
 assign la_data_out[20] = net258;
 assign la_data_out[21] = net259;
 assign la_data_out[22] = net260;
 assign la_data_out[23] = net261;
 assign la_data_out[24] = net262;
 assign la_data_out[25] = net263;
 assign la_data_out[26] = net264;
 assign la_data_out[27] = net265;
 assign la_data_out[28] = net266;
 assign la_data_out[29] = net267;
 assign la_data_out[2] = net240;
 assign la_data_out[30] = net268;
 assign la_data_out[31] = net269;
 assign la_data_out[32] = net270;
 assign la_data_out[33] = net271;
 assign la_data_out[34] = net272;
 assign la_data_out[35] = net273;
 assign la_data_out[36] = net274;
 assign la_data_out[37] = net275;
 assign la_data_out[38] = net276;
 assign la_data_out[39] = net277;
 assign la_data_out[3] = net241;
 assign la_data_out[40] = net278;
 assign la_data_out[41] = net279;
 assign la_data_out[42] = net280;
 assign la_data_out[43] = net281;
 assign la_data_out[44] = net282;
 assign la_data_out[45] = net283;
 assign la_data_out[46] = net284;
 assign la_data_out[47] = net285;
 assign la_data_out[48] = net286;
 assign la_data_out[49] = net287;
 assign la_data_out[4] = net242;
 assign la_data_out[50] = net288;
 assign la_data_out[51] = net289;
 assign la_data_out[52] = net290;
 assign la_data_out[53] = net291;
 assign la_data_out[54] = net292;
 assign la_data_out[55] = net293;
 assign la_data_out[56] = net294;
 assign la_data_out[57] = net295;
 assign la_data_out[58] = net296;
 assign la_data_out[59] = net297;
 assign la_data_out[5] = net243;
 assign la_data_out[60] = net298;
 assign la_data_out[61] = net299;
 assign la_data_out[62] = net300;
 assign la_data_out[63] = net301;
 assign la_data_out[64] = net302;
 assign la_data_out[65] = net303;
 assign la_data_out[66] = net304;
 assign la_data_out[67] = net305;
 assign la_data_out[68] = net306;
 assign la_data_out[69] = net307;
 assign la_data_out[6] = net244;
 assign la_data_out[70] = net308;
 assign la_data_out[71] = net309;
 assign la_data_out[72] = net310;
 assign la_data_out[73] = net311;
 assign la_data_out[74] = net312;
 assign la_data_out[75] = net313;
 assign la_data_out[76] = net314;
 assign la_data_out[77] = net315;
 assign la_data_out[78] = net316;
 assign la_data_out[79] = net317;
 assign la_data_out[7] = net245;
 assign la_data_out[80] = net318;
 assign la_data_out[81] = net319;
 assign la_data_out[82] = net320;
 assign la_data_out[83] = net321;
 assign la_data_out[84] = net322;
 assign la_data_out[85] = net323;
 assign la_data_out[86] = net324;
 assign la_data_out[87] = net325;
 assign la_data_out[88] = net326;
 assign la_data_out[89] = net327;
 assign la_data_out[8] = net246;
 assign la_data_out[90] = net328;
 assign la_data_out[91] = net329;
 assign la_data_out[92] = net330;
 assign la_data_out[93] = net331;
 assign la_data_out[94] = net332;
 assign la_data_out[95] = net333;
 assign la_data_out[96] = net334;
 assign la_data_out[97] = net335;
 assign la_data_out[98] = net336;
 assign la_data_out[99] = net337;
 assign la_data_out[9] = net247;
 assign m_io_oeb[26] = net414;
 assign m_io_oeb[27] = net415;
 assign m_io_oeb[28] = net368;
 assign m_io_oeb[29] = net369;
 assign m_io_oeb[30] = net416;
 assign m_io_oeb[31] = net417;
 assign m_io_oeb[32] = net418;
 assign m_io_oeb[33] = net419;
 assign m_io_oeb[34] = net420;
 assign m_io_oeb[35] = net421;
 assign m_io_oeb[36] = net370;
 assign m_io_oeb[37] = net371;
 assign m_io_oeb[8] = net366;
 assign m_io_oeb[9] = net367;
 assign m_io_out[26] = net372;
 assign m_io_out[27] = net373;
 assign m_io_out[30] = net374;
 assign m_io_out[31] = net375;
 assign m_io_out[32] = net376;
 assign m_io_out[33] = net377;
 assign m_io_out[34] = net378;
 assign m_io_out[35] = net379;
 assign m_io_out[37] = net422;
 assign mgt_wb_ack_o = net380;
 assign mgt_wb_dat_o[0] = net381;
 assign mgt_wb_dat_o[10] = net391;
 assign mgt_wb_dat_o[11] = net392;
 assign mgt_wb_dat_o[12] = net393;
 assign mgt_wb_dat_o[13] = net394;
 assign mgt_wb_dat_o[14] = net395;
 assign mgt_wb_dat_o[15] = net396;
 assign mgt_wb_dat_o[16] = net397;
 assign mgt_wb_dat_o[17] = net398;
 assign mgt_wb_dat_o[18] = net399;
 assign mgt_wb_dat_o[19] = net400;
 assign mgt_wb_dat_o[1] = net382;
 assign mgt_wb_dat_o[20] = net401;
 assign mgt_wb_dat_o[21] = net402;
 assign mgt_wb_dat_o[22] = net403;
 assign mgt_wb_dat_o[23] = net404;
 assign mgt_wb_dat_o[24] = net405;
 assign mgt_wb_dat_o[25] = net406;
 assign mgt_wb_dat_o[26] = net407;
 assign mgt_wb_dat_o[27] = net408;
 assign mgt_wb_dat_o[28] = net409;
 assign mgt_wb_dat_o[29] = net410;
 assign mgt_wb_dat_o[2] = net383;
 assign mgt_wb_dat_o[30] = net411;
 assign mgt_wb_dat_o[31] = net412;
 assign mgt_wb_dat_o[3] = net384;
 assign mgt_wb_dat_o[4] = net385;
 assign mgt_wb_dat_o[5] = net386;
 assign mgt_wb_dat_o[6] = net387;
 assign mgt_wb_dat_o[7] = net388;
 assign mgt_wb_dat_o[8] = net389;
 assign mgt_wb_dat_o[9] = net390;
endmodule

