magic
tech sky130A
magscale 1 2
timestamp 1672399398
<< nwell >>
rect 1066 77509 58918 77830
rect 1066 76421 58918 76987
rect 1066 75333 58918 75899
rect 1066 74245 58918 74811
rect 1066 73157 58918 73723
rect 1066 72069 58918 72635
rect 1066 70981 58918 71547
rect 1066 69893 58918 70459
rect 1066 68805 58918 69371
rect 1066 67717 58918 68283
rect 1066 66629 58918 67195
rect 1066 65541 58918 66107
rect 1066 64453 58918 65019
rect 1066 63365 58918 63931
rect 1066 62277 58918 62843
rect 1066 61189 58918 61755
rect 1066 60101 58918 60667
rect 1066 59013 58918 59579
rect 1066 57925 58918 58491
rect 1066 56837 58918 57403
rect 1066 55749 58918 56315
rect 1066 54661 58918 55227
rect 1066 53573 58918 54139
rect 1066 52485 58918 53051
rect 1066 51397 58918 51963
rect 1066 50309 58918 50875
rect 1066 49221 58918 49787
rect 1066 48133 58918 48699
rect 1066 47045 58918 47611
rect 1066 45957 58918 46523
rect 1066 44869 58918 45435
rect 1066 43781 58918 44347
rect 1066 42693 58918 43259
rect 1066 41605 58918 42171
rect 1066 40517 58918 41083
rect 1066 39429 58918 39995
rect 1066 38341 58918 38907
rect 1066 37253 58918 37819
rect 1066 36165 58918 36731
rect 1066 35077 58918 35643
rect 1066 33989 58918 34555
rect 1066 32901 58918 33467
rect 1066 31813 58918 32379
rect 1066 30725 58918 31291
rect 1066 29637 58918 30203
rect 1066 28549 58918 29115
rect 1066 27461 58918 28027
rect 1066 26373 58918 26939
rect 1066 25285 58918 25851
rect 1066 24197 58918 24763
rect 1066 23109 58918 23675
rect 1066 22021 58918 22587
rect 1066 20933 58918 21499
rect 1066 19845 58918 20411
rect 1066 18757 58918 19323
rect 1066 17669 58918 18235
rect 1066 16581 58918 17147
rect 1066 15493 58918 16059
rect 1066 14405 58918 14971
rect 1066 13317 58918 13883
rect 1066 12229 58918 12795
rect 1066 11141 58918 11707
rect 1066 10053 58918 10619
rect 1066 8965 58918 9531
rect 1066 7877 58918 8443
rect 1066 6789 58918 7355
rect 1066 5701 58918 6267
rect 1066 4613 58918 5179
rect 1066 3525 58918 4091
rect 1066 2437 58918 3003
<< obsli1 >>
rect 1104 2159 58880 77809
<< obsm1 >>
rect 1104 1844 58880 78940
<< metal2 >>
rect 2042 79200 2098 80000
rect 2134 79200 2190 80000
rect 2226 79200 2282 80000
rect 2318 79200 2374 80000
rect 2410 79200 2466 80000
rect 2502 79200 2558 80000
rect 2594 79200 2650 80000
rect 2686 79200 2742 80000
rect 2778 79200 2834 80000
rect 2870 79200 2926 80000
rect 2962 79200 3018 80000
rect 3054 79200 3110 80000
rect 3146 79200 3202 80000
rect 3238 79200 3294 80000
rect 3330 79200 3386 80000
rect 3422 79200 3478 80000
rect 3514 79200 3570 80000
rect 3606 79200 3662 80000
rect 3698 79200 3754 80000
rect 3790 79200 3846 80000
rect 3882 79200 3938 80000
rect 3974 79200 4030 80000
rect 4066 79200 4122 80000
rect 4158 79200 4214 80000
rect 4250 79200 4306 80000
rect 4342 79200 4398 80000
rect 4434 79200 4490 80000
rect 4526 79200 4582 80000
rect 4618 79200 4674 80000
rect 4710 79200 4766 80000
rect 4802 79200 4858 80000
rect 4894 79200 4950 80000
rect 4986 79200 5042 80000
rect 5078 79200 5134 80000
rect 5170 79200 5226 80000
rect 5262 79200 5318 80000
rect 5354 79200 5410 80000
rect 5446 79200 5502 80000
rect 5538 79200 5594 80000
rect 5630 79200 5686 80000
rect 5722 79200 5778 80000
rect 5814 79200 5870 80000
rect 5906 79200 5962 80000
rect 5998 79200 6054 80000
rect 6090 79200 6146 80000
rect 6182 79200 6238 80000
rect 6274 79200 6330 80000
rect 6366 79200 6422 80000
rect 6458 79200 6514 80000
rect 6550 79200 6606 80000
rect 6642 79200 6698 80000
rect 6734 79200 6790 80000
rect 6826 79200 6882 80000
rect 6918 79200 6974 80000
rect 7010 79200 7066 80000
rect 7102 79200 7158 80000
rect 7194 79200 7250 80000
rect 7286 79200 7342 80000
rect 7378 79200 7434 80000
rect 7470 79200 7526 80000
rect 7562 79200 7618 80000
rect 7654 79200 7710 80000
rect 7746 79200 7802 80000
rect 7838 79200 7894 80000
rect 7930 79200 7986 80000
rect 8022 79200 8078 80000
rect 8114 79200 8170 80000
rect 8206 79200 8262 80000
rect 8298 79200 8354 80000
rect 8390 79200 8446 80000
rect 8482 79200 8538 80000
rect 8574 79200 8630 80000
rect 8666 79200 8722 80000
rect 8758 79200 8814 80000
rect 8850 79200 8906 80000
rect 8942 79200 8998 80000
rect 9034 79200 9090 80000
rect 9126 79200 9182 80000
rect 9218 79200 9274 80000
rect 9310 79200 9366 80000
rect 9402 79200 9458 80000
rect 9494 79200 9550 80000
rect 9586 79200 9642 80000
rect 9678 79200 9734 80000
rect 9770 79200 9826 80000
rect 9862 79200 9918 80000
rect 9954 79200 10010 80000
rect 10046 79200 10102 80000
rect 10138 79200 10194 80000
rect 10230 79200 10286 80000
rect 10322 79200 10378 80000
rect 10414 79200 10470 80000
rect 10506 79200 10562 80000
rect 10598 79200 10654 80000
rect 10690 79200 10746 80000
rect 10782 79200 10838 80000
rect 10874 79200 10930 80000
rect 10966 79200 11022 80000
rect 11058 79200 11114 80000
rect 11150 79200 11206 80000
rect 11242 79200 11298 80000
rect 11334 79200 11390 80000
rect 11426 79200 11482 80000
rect 11518 79200 11574 80000
rect 11610 79200 11666 80000
rect 11702 79200 11758 80000
rect 11794 79200 11850 80000
rect 11886 79200 11942 80000
rect 11978 79200 12034 80000
rect 12070 79200 12126 80000
rect 12162 79200 12218 80000
rect 12254 79200 12310 80000
rect 12346 79200 12402 80000
rect 12438 79200 12494 80000
rect 12530 79200 12586 80000
rect 12622 79200 12678 80000
rect 12714 79200 12770 80000
rect 12806 79200 12862 80000
rect 12898 79200 12954 80000
rect 12990 79200 13046 80000
rect 13082 79200 13138 80000
rect 13174 79200 13230 80000
rect 13266 79200 13322 80000
rect 13358 79200 13414 80000
rect 13450 79200 13506 80000
rect 13542 79200 13598 80000
rect 13634 79200 13690 80000
rect 13726 79200 13782 80000
rect 13818 79200 13874 80000
rect 13910 79200 13966 80000
rect 14002 79200 14058 80000
rect 14094 79200 14150 80000
rect 14186 79200 14242 80000
rect 14278 79200 14334 80000
rect 14370 79200 14426 80000
rect 14462 79200 14518 80000
rect 14554 79200 14610 80000
rect 14646 79200 14702 80000
rect 14738 79200 14794 80000
rect 14830 79200 14886 80000
rect 14922 79200 14978 80000
rect 15014 79200 15070 80000
rect 15106 79200 15162 80000
rect 15198 79200 15254 80000
rect 15290 79200 15346 80000
rect 15382 79200 15438 80000
rect 15474 79200 15530 80000
rect 15566 79200 15622 80000
rect 15658 79200 15714 80000
rect 15750 79200 15806 80000
rect 15842 79200 15898 80000
rect 15934 79200 15990 80000
rect 16026 79200 16082 80000
rect 16118 79200 16174 80000
rect 16210 79200 16266 80000
rect 16302 79200 16358 80000
rect 16394 79200 16450 80000
rect 16486 79200 16542 80000
rect 16578 79200 16634 80000
rect 16670 79200 16726 80000
rect 16762 79200 16818 80000
rect 16854 79200 16910 80000
rect 16946 79200 17002 80000
rect 17038 79200 17094 80000
rect 17130 79200 17186 80000
rect 17222 79200 17278 80000
rect 17314 79200 17370 80000
rect 17406 79200 17462 80000
rect 17498 79200 17554 80000
rect 17590 79200 17646 80000
rect 17682 79200 17738 80000
rect 17774 79200 17830 80000
rect 17866 79200 17922 80000
rect 17958 79200 18014 80000
rect 18050 79200 18106 80000
rect 18142 79200 18198 80000
rect 18234 79200 18290 80000
rect 18326 79200 18382 80000
rect 18418 79200 18474 80000
rect 18510 79200 18566 80000
rect 18602 79200 18658 80000
rect 18694 79200 18750 80000
rect 18786 79200 18842 80000
rect 18878 79200 18934 80000
rect 18970 79200 19026 80000
rect 19062 79200 19118 80000
rect 19154 79200 19210 80000
rect 19246 79200 19302 80000
rect 19338 79200 19394 80000
rect 19430 79200 19486 80000
rect 19522 79200 19578 80000
rect 19614 79200 19670 80000
rect 19706 79200 19762 80000
rect 19798 79200 19854 80000
rect 19890 79200 19946 80000
rect 19982 79200 20038 80000
rect 20074 79200 20130 80000
rect 20166 79200 20222 80000
rect 20258 79200 20314 80000
rect 20350 79200 20406 80000
rect 20442 79200 20498 80000
rect 20534 79200 20590 80000
rect 20626 79200 20682 80000
rect 20718 79200 20774 80000
rect 20810 79200 20866 80000
rect 20902 79200 20958 80000
rect 20994 79200 21050 80000
rect 21086 79200 21142 80000
rect 21178 79200 21234 80000
rect 21270 79200 21326 80000
rect 21362 79200 21418 80000
rect 21454 79200 21510 80000
rect 21546 79200 21602 80000
rect 21638 79200 21694 80000
rect 21730 79200 21786 80000
rect 21822 79200 21878 80000
rect 21914 79200 21970 80000
rect 22006 79200 22062 80000
rect 22098 79200 22154 80000
rect 22190 79200 22246 80000
rect 22282 79200 22338 80000
rect 22374 79200 22430 80000
rect 22466 79200 22522 80000
rect 22558 79200 22614 80000
rect 22650 79200 22706 80000
rect 22742 79200 22798 80000
rect 22834 79200 22890 80000
rect 22926 79200 22982 80000
rect 23018 79200 23074 80000
rect 23110 79200 23166 80000
rect 23202 79200 23258 80000
rect 23294 79200 23350 80000
rect 23386 79200 23442 80000
rect 23478 79200 23534 80000
rect 23570 79200 23626 80000
rect 23662 79200 23718 80000
rect 23754 79200 23810 80000
rect 23846 79200 23902 80000
rect 23938 79200 23994 80000
rect 24030 79200 24086 80000
rect 24122 79200 24178 80000
rect 24214 79200 24270 80000
rect 24306 79200 24362 80000
rect 24398 79200 24454 80000
rect 24490 79200 24546 80000
rect 24582 79200 24638 80000
rect 24674 79200 24730 80000
rect 24766 79200 24822 80000
rect 24858 79200 24914 80000
rect 24950 79200 25006 80000
rect 25042 79200 25098 80000
rect 25134 79200 25190 80000
rect 25226 79200 25282 80000
rect 25318 79200 25374 80000
rect 25410 79200 25466 80000
rect 25502 79200 25558 80000
rect 25594 79200 25650 80000
rect 25686 79200 25742 80000
rect 25778 79200 25834 80000
rect 25870 79200 25926 80000
rect 25962 79200 26018 80000
rect 26054 79200 26110 80000
rect 26146 79200 26202 80000
rect 26238 79200 26294 80000
rect 26330 79200 26386 80000
rect 26422 79200 26478 80000
rect 26514 79200 26570 80000
rect 26606 79200 26662 80000
rect 26698 79200 26754 80000
rect 26790 79200 26846 80000
rect 26882 79200 26938 80000
rect 26974 79200 27030 80000
rect 27066 79200 27122 80000
rect 27158 79200 27214 80000
rect 27250 79200 27306 80000
rect 27342 79200 27398 80000
rect 27434 79200 27490 80000
rect 27526 79200 27582 80000
rect 27618 79200 27674 80000
rect 27710 79200 27766 80000
rect 27802 79200 27858 80000
rect 27894 79200 27950 80000
rect 27986 79200 28042 80000
rect 28078 79200 28134 80000
rect 28170 79200 28226 80000
rect 28262 79200 28318 80000
rect 28354 79200 28410 80000
rect 28446 79200 28502 80000
rect 28538 79200 28594 80000
rect 28630 79200 28686 80000
rect 28722 79200 28778 80000
rect 28814 79200 28870 80000
rect 28906 79200 28962 80000
rect 28998 79200 29054 80000
rect 29090 79200 29146 80000
rect 29182 79200 29238 80000
rect 29274 79200 29330 80000
rect 29366 79200 29422 80000
rect 29458 79200 29514 80000
rect 29550 79200 29606 80000
rect 29642 79200 29698 80000
rect 29734 79200 29790 80000
rect 29826 79200 29882 80000
rect 29918 79200 29974 80000
rect 30010 79200 30066 80000
rect 30102 79200 30158 80000
rect 30194 79200 30250 80000
rect 30286 79200 30342 80000
rect 30378 79200 30434 80000
rect 30470 79200 30526 80000
rect 30562 79200 30618 80000
rect 30654 79200 30710 80000
rect 30746 79200 30802 80000
rect 30838 79200 30894 80000
rect 30930 79200 30986 80000
rect 31022 79200 31078 80000
rect 31114 79200 31170 80000
rect 31206 79200 31262 80000
rect 31298 79200 31354 80000
rect 31390 79200 31446 80000
rect 31482 79200 31538 80000
rect 31574 79200 31630 80000
rect 31666 79200 31722 80000
rect 31758 79200 31814 80000
rect 31850 79200 31906 80000
rect 31942 79200 31998 80000
rect 32034 79200 32090 80000
rect 32126 79200 32182 80000
rect 32218 79200 32274 80000
rect 32310 79200 32366 80000
rect 32402 79200 32458 80000
rect 32494 79200 32550 80000
rect 32586 79200 32642 80000
rect 32678 79200 32734 80000
rect 32770 79200 32826 80000
rect 32862 79200 32918 80000
rect 32954 79200 33010 80000
rect 33046 79200 33102 80000
rect 33138 79200 33194 80000
rect 33230 79200 33286 80000
rect 33322 79200 33378 80000
rect 33414 79200 33470 80000
rect 33506 79200 33562 80000
rect 33598 79200 33654 80000
rect 33690 79200 33746 80000
rect 33782 79200 33838 80000
rect 33874 79200 33930 80000
rect 33966 79200 34022 80000
rect 34058 79200 34114 80000
rect 34150 79200 34206 80000
rect 34242 79200 34298 80000
rect 34334 79200 34390 80000
rect 34426 79200 34482 80000
rect 34518 79200 34574 80000
rect 34610 79200 34666 80000
rect 34702 79200 34758 80000
rect 34794 79200 34850 80000
rect 34886 79200 34942 80000
rect 34978 79200 35034 80000
rect 35070 79200 35126 80000
rect 35162 79200 35218 80000
rect 35254 79200 35310 80000
rect 35346 79200 35402 80000
rect 35438 79200 35494 80000
rect 35530 79200 35586 80000
rect 35622 79200 35678 80000
rect 35714 79200 35770 80000
rect 35806 79200 35862 80000
rect 35898 79200 35954 80000
rect 35990 79200 36046 80000
rect 36082 79200 36138 80000
rect 36174 79200 36230 80000
rect 36266 79200 36322 80000
rect 36358 79200 36414 80000
rect 36450 79200 36506 80000
rect 36542 79200 36598 80000
rect 36634 79200 36690 80000
rect 36726 79200 36782 80000
rect 36818 79200 36874 80000
rect 36910 79200 36966 80000
rect 37002 79200 37058 80000
rect 37094 79200 37150 80000
rect 37186 79200 37242 80000
rect 37278 79200 37334 80000
rect 37370 79200 37426 80000
rect 37462 79200 37518 80000
rect 37554 79200 37610 80000
rect 37646 79200 37702 80000
rect 37738 79200 37794 80000
rect 37830 79200 37886 80000
rect 37922 79200 37978 80000
rect 38014 79200 38070 80000
rect 38106 79200 38162 80000
rect 38198 79200 38254 80000
rect 38290 79200 38346 80000
rect 38382 79200 38438 80000
rect 38474 79200 38530 80000
rect 38566 79200 38622 80000
rect 38658 79200 38714 80000
rect 38750 79200 38806 80000
rect 38842 79200 38898 80000
rect 38934 79200 38990 80000
rect 39026 79200 39082 80000
rect 39118 79200 39174 80000
rect 39210 79200 39266 80000
rect 39302 79200 39358 80000
rect 39394 79200 39450 80000
rect 39486 79200 39542 80000
rect 39578 79200 39634 80000
rect 39670 79200 39726 80000
rect 39762 79200 39818 80000
rect 39854 79200 39910 80000
rect 39946 79200 40002 80000
rect 40038 79200 40094 80000
rect 40130 79200 40186 80000
rect 40222 79200 40278 80000
rect 40314 79200 40370 80000
rect 40406 79200 40462 80000
rect 40498 79200 40554 80000
rect 40590 79200 40646 80000
rect 40682 79200 40738 80000
rect 40774 79200 40830 80000
rect 40866 79200 40922 80000
rect 40958 79200 41014 80000
rect 41050 79200 41106 80000
rect 41142 79200 41198 80000
rect 41234 79200 41290 80000
rect 41326 79200 41382 80000
rect 41418 79200 41474 80000
rect 41510 79200 41566 80000
rect 41602 79200 41658 80000
rect 41694 79200 41750 80000
rect 41786 79200 41842 80000
rect 41878 79200 41934 80000
rect 41970 79200 42026 80000
rect 42062 79200 42118 80000
rect 42154 79200 42210 80000
rect 42246 79200 42302 80000
rect 42338 79200 42394 80000
rect 42430 79200 42486 80000
rect 42522 79200 42578 80000
rect 42614 79200 42670 80000
rect 42706 79200 42762 80000
rect 42798 79200 42854 80000
rect 42890 79200 42946 80000
rect 42982 79200 43038 80000
rect 43074 79200 43130 80000
rect 43166 79200 43222 80000
rect 43258 79200 43314 80000
rect 43350 79200 43406 80000
rect 43442 79200 43498 80000
rect 43534 79200 43590 80000
rect 43626 79200 43682 80000
rect 43718 79200 43774 80000
rect 43810 79200 43866 80000
rect 43902 79200 43958 80000
rect 43994 79200 44050 80000
rect 44086 79200 44142 80000
rect 44178 79200 44234 80000
rect 44270 79200 44326 80000
rect 44362 79200 44418 80000
rect 44454 79200 44510 80000
rect 44546 79200 44602 80000
rect 44638 79200 44694 80000
rect 44730 79200 44786 80000
rect 44822 79200 44878 80000
rect 44914 79200 44970 80000
rect 45006 79200 45062 80000
rect 45098 79200 45154 80000
rect 45190 79200 45246 80000
rect 45282 79200 45338 80000
rect 45374 79200 45430 80000
rect 45466 79200 45522 80000
rect 45558 79200 45614 80000
rect 45650 79200 45706 80000
rect 45742 79200 45798 80000
rect 45834 79200 45890 80000
rect 45926 79200 45982 80000
rect 46018 79200 46074 80000
rect 46110 79200 46166 80000
rect 46202 79200 46258 80000
rect 46294 79200 46350 80000
rect 46386 79200 46442 80000
rect 46478 79200 46534 80000
rect 46570 79200 46626 80000
rect 46662 79200 46718 80000
rect 46754 79200 46810 80000
rect 46846 79200 46902 80000
rect 46938 79200 46994 80000
rect 47030 79200 47086 80000
rect 47122 79200 47178 80000
rect 47214 79200 47270 80000
rect 47306 79200 47362 80000
rect 47398 79200 47454 80000
rect 47490 79200 47546 80000
rect 47582 79200 47638 80000
rect 47674 79200 47730 80000
rect 47766 79200 47822 80000
rect 47858 79200 47914 80000
rect 47950 79200 48006 80000
rect 48042 79200 48098 80000
rect 48134 79200 48190 80000
rect 48226 79200 48282 80000
rect 48318 79200 48374 80000
rect 48410 79200 48466 80000
rect 48502 79200 48558 80000
rect 48594 79200 48650 80000
rect 48686 79200 48742 80000
rect 48778 79200 48834 80000
rect 48870 79200 48926 80000
rect 48962 79200 49018 80000
rect 49054 79200 49110 80000
rect 49146 79200 49202 80000
rect 49238 79200 49294 80000
rect 49330 79200 49386 80000
rect 49422 79200 49478 80000
rect 49514 79200 49570 80000
rect 49606 79200 49662 80000
rect 49698 79200 49754 80000
rect 49790 79200 49846 80000
rect 49882 79200 49938 80000
rect 49974 79200 50030 80000
rect 50066 79200 50122 80000
rect 50158 79200 50214 80000
rect 50250 79200 50306 80000
rect 50342 79200 50398 80000
rect 50434 79200 50490 80000
rect 50526 79200 50582 80000
rect 50618 79200 50674 80000
rect 50710 79200 50766 80000
rect 50802 79200 50858 80000
rect 50894 79200 50950 80000
rect 50986 79200 51042 80000
rect 51078 79200 51134 80000
rect 51170 79200 51226 80000
rect 51262 79200 51318 80000
rect 51354 79200 51410 80000
rect 51446 79200 51502 80000
rect 51538 79200 51594 80000
rect 51630 79200 51686 80000
rect 51722 79200 51778 80000
rect 51814 79200 51870 80000
rect 51906 79200 51962 80000
rect 51998 79200 52054 80000
rect 52090 79200 52146 80000
rect 52182 79200 52238 80000
rect 52274 79200 52330 80000
rect 52366 79200 52422 80000
rect 52458 79200 52514 80000
rect 52550 79200 52606 80000
rect 52642 79200 52698 80000
rect 52734 79200 52790 80000
rect 52826 79200 52882 80000
rect 52918 79200 52974 80000
rect 53010 79200 53066 80000
rect 53102 79200 53158 80000
rect 53194 79200 53250 80000
rect 53286 79200 53342 80000
rect 53378 79200 53434 80000
rect 53470 79200 53526 80000
rect 53562 79200 53618 80000
rect 53654 79200 53710 80000
rect 53746 79200 53802 80000
rect 53838 79200 53894 80000
rect 53930 79200 53986 80000
rect 54022 79200 54078 80000
rect 54114 79200 54170 80000
rect 54206 79200 54262 80000
rect 54298 79200 54354 80000
rect 54390 79200 54446 80000
rect 54482 79200 54538 80000
rect 54574 79200 54630 80000
rect 54666 79200 54722 80000
rect 54758 79200 54814 80000
rect 54850 79200 54906 80000
rect 54942 79200 54998 80000
rect 55034 79200 55090 80000
rect 55126 79200 55182 80000
rect 55218 79200 55274 80000
rect 55310 79200 55366 80000
rect 55402 79200 55458 80000
rect 55494 79200 55550 80000
rect 55586 79200 55642 80000
rect 55678 79200 55734 80000
rect 55770 79200 55826 80000
rect 55862 79200 55918 80000
rect 55954 79200 56010 80000
rect 56046 79200 56102 80000
rect 56138 79200 56194 80000
rect 56230 79200 56286 80000
rect 56322 79200 56378 80000
rect 56414 79200 56470 80000
rect 56506 79200 56562 80000
rect 56598 79200 56654 80000
rect 56690 79200 56746 80000
rect 56782 79200 56838 80000
rect 56874 79200 56930 80000
rect 56966 79200 57022 80000
rect 57058 79200 57114 80000
rect 57150 79200 57206 80000
rect 57242 79200 57298 80000
rect 57334 79200 57390 80000
rect 57426 79200 57482 80000
rect 57518 79200 57574 80000
rect 57610 79200 57666 80000
rect 57702 79200 57758 80000
rect 57794 79200 57850 80000
rect 57886 79200 57942 80000
rect 1398 0 1454 800
rect 2226 0 2282 800
rect 3054 0 3110 800
rect 3882 0 3938 800
rect 4710 0 4766 800
rect 5538 0 5594 800
rect 6366 0 6422 800
rect 7194 0 7250 800
rect 8022 0 8078 800
rect 8850 0 8906 800
rect 9678 0 9734 800
rect 10506 0 10562 800
rect 11334 0 11390 800
rect 12162 0 12218 800
rect 12990 0 13046 800
rect 13818 0 13874 800
rect 14646 0 14702 800
rect 15474 0 15530 800
rect 16302 0 16358 800
rect 17130 0 17186 800
rect 17958 0 18014 800
rect 18786 0 18842 800
rect 19614 0 19670 800
rect 20442 0 20498 800
rect 21270 0 21326 800
rect 22098 0 22154 800
rect 22926 0 22982 800
rect 23754 0 23810 800
rect 24582 0 24638 800
rect 25410 0 25466 800
rect 26238 0 26294 800
rect 27066 0 27122 800
rect 27894 0 27950 800
rect 28722 0 28778 800
rect 29550 0 29606 800
rect 30378 0 30434 800
rect 31206 0 31262 800
rect 32034 0 32090 800
rect 32862 0 32918 800
rect 33690 0 33746 800
rect 34518 0 34574 800
rect 35346 0 35402 800
rect 36174 0 36230 800
rect 37002 0 37058 800
rect 37830 0 37886 800
rect 38658 0 38714 800
rect 39486 0 39542 800
rect 40314 0 40370 800
rect 41142 0 41198 800
rect 41970 0 42026 800
rect 42798 0 42854 800
rect 43626 0 43682 800
rect 44454 0 44510 800
rect 45282 0 45338 800
rect 46110 0 46166 800
rect 46938 0 46994 800
rect 47766 0 47822 800
rect 48594 0 48650 800
rect 49422 0 49478 800
rect 50250 0 50306 800
rect 51078 0 51134 800
rect 51906 0 51962 800
rect 52734 0 52790 800
rect 53562 0 53618 800
rect 54390 0 54446 800
rect 55218 0 55274 800
rect 56046 0 56102 800
rect 56874 0 56930 800
rect 57702 0 57758 800
rect 58530 0 58586 800
<< obsm2 >>
rect 1400 79144 1986 79200
rect 57998 79144 58676 79200
rect 1400 856 58676 79144
rect 1510 734 2170 856
rect 2338 734 2998 856
rect 3166 734 3826 856
rect 3994 734 4654 856
rect 4822 734 5482 856
rect 5650 734 6310 856
rect 6478 734 7138 856
rect 7306 734 7966 856
rect 8134 734 8794 856
rect 8962 734 9622 856
rect 9790 734 10450 856
rect 10618 734 11278 856
rect 11446 734 12106 856
rect 12274 734 12934 856
rect 13102 734 13762 856
rect 13930 734 14590 856
rect 14758 734 15418 856
rect 15586 734 16246 856
rect 16414 734 17074 856
rect 17242 734 17902 856
rect 18070 734 18730 856
rect 18898 734 19558 856
rect 19726 734 20386 856
rect 20554 734 21214 856
rect 21382 734 22042 856
rect 22210 734 22870 856
rect 23038 734 23698 856
rect 23866 734 24526 856
rect 24694 734 25354 856
rect 25522 734 26182 856
rect 26350 734 27010 856
rect 27178 734 27838 856
rect 28006 734 28666 856
rect 28834 734 29494 856
rect 29662 734 30322 856
rect 30490 734 31150 856
rect 31318 734 31978 856
rect 32146 734 32806 856
rect 32974 734 33634 856
rect 33802 734 34462 856
rect 34630 734 35290 856
rect 35458 734 36118 856
rect 36286 734 36946 856
rect 37114 734 37774 856
rect 37942 734 38602 856
rect 38770 734 39430 856
rect 39598 734 40258 856
rect 40426 734 41086 856
rect 41254 734 41914 856
rect 42082 734 42742 856
rect 42910 734 43570 856
rect 43738 734 44398 856
rect 44566 734 45226 856
rect 45394 734 46054 856
rect 46222 734 46882 856
rect 47050 734 47710 856
rect 47878 734 48538 856
rect 48706 734 49366 856
rect 49534 734 50194 856
rect 50362 734 51022 856
rect 51190 734 51850 856
rect 52018 734 52678 856
rect 52846 734 53506 856
rect 53674 734 54334 856
rect 54502 734 55162 856
rect 55330 734 55990 856
rect 56158 734 56818 856
rect 56986 734 57646 856
rect 57814 734 58474 856
rect 58642 734 58676 856
<< metal3 >>
rect 59200 72496 60000 72616
rect 59200 71952 60000 72072
rect 59200 71408 60000 71528
rect 59200 70864 60000 70984
rect 59200 70320 60000 70440
rect 59200 69776 60000 69896
rect 59200 69232 60000 69352
rect 59200 68688 60000 68808
rect 59200 68144 60000 68264
rect 59200 67600 60000 67720
rect 59200 67056 60000 67176
rect 59200 66512 60000 66632
rect 59200 65968 60000 66088
rect 59200 65424 60000 65544
rect 59200 64880 60000 65000
rect 59200 64336 60000 64456
rect 59200 63792 60000 63912
rect 59200 63248 60000 63368
rect 59200 62704 60000 62824
rect 59200 62160 60000 62280
rect 59200 61616 60000 61736
rect 59200 61072 60000 61192
rect 59200 60528 60000 60648
rect 59200 59984 60000 60104
rect 59200 59440 60000 59560
rect 59200 58896 60000 59016
rect 59200 58352 60000 58472
rect 59200 57808 60000 57928
rect 59200 57264 60000 57384
rect 59200 56720 60000 56840
rect 59200 56176 60000 56296
rect 59200 55632 60000 55752
rect 59200 55088 60000 55208
rect 59200 54544 60000 54664
rect 59200 54000 60000 54120
rect 59200 53456 60000 53576
rect 59200 52912 60000 53032
rect 59200 52368 60000 52488
rect 59200 51824 60000 51944
rect 59200 51280 60000 51400
rect 59200 50736 60000 50856
rect 59200 50192 60000 50312
rect 59200 49648 60000 49768
rect 59200 49104 60000 49224
rect 59200 48560 60000 48680
rect 59200 48016 60000 48136
rect 59200 47472 60000 47592
rect 59200 46928 60000 47048
rect 59200 46384 60000 46504
rect 59200 45840 60000 45960
rect 59200 45296 60000 45416
rect 59200 44752 60000 44872
rect 59200 44208 60000 44328
rect 59200 43664 60000 43784
rect 59200 43120 60000 43240
rect 59200 42576 60000 42696
rect 59200 42032 60000 42152
rect 59200 41488 60000 41608
rect 59200 40944 60000 41064
rect 59200 40400 60000 40520
rect 59200 39856 60000 39976
rect 59200 39312 60000 39432
rect 59200 38768 60000 38888
rect 59200 38224 60000 38344
rect 59200 37680 60000 37800
rect 59200 37136 60000 37256
rect 59200 36592 60000 36712
rect 59200 36048 60000 36168
rect 59200 35504 60000 35624
rect 59200 34960 60000 35080
rect 59200 34416 60000 34536
rect 59200 33872 60000 33992
rect 59200 33328 60000 33448
rect 59200 32784 60000 32904
rect 59200 32240 60000 32360
rect 59200 31696 60000 31816
rect 59200 31152 60000 31272
rect 59200 30608 60000 30728
rect 59200 30064 60000 30184
rect 59200 29520 60000 29640
rect 59200 28976 60000 29096
rect 59200 28432 60000 28552
rect 59200 27888 60000 28008
rect 59200 27344 60000 27464
rect 59200 26800 60000 26920
rect 59200 26256 60000 26376
rect 59200 25712 60000 25832
rect 59200 25168 60000 25288
rect 59200 24624 60000 24744
rect 59200 24080 60000 24200
rect 59200 23536 60000 23656
rect 59200 22992 60000 23112
rect 59200 22448 60000 22568
rect 59200 21904 60000 22024
rect 59200 21360 60000 21480
rect 59200 20816 60000 20936
rect 59200 20272 60000 20392
rect 59200 19728 60000 19848
rect 59200 19184 60000 19304
rect 59200 18640 60000 18760
rect 59200 18096 60000 18216
rect 59200 17552 60000 17672
rect 59200 17008 60000 17128
rect 59200 16464 60000 16584
rect 59200 15920 60000 16040
rect 59200 15376 60000 15496
rect 59200 14832 60000 14952
rect 59200 14288 60000 14408
rect 59200 13744 60000 13864
rect 59200 13200 60000 13320
rect 59200 12656 60000 12776
rect 59200 12112 60000 12232
rect 59200 11568 60000 11688
rect 59200 11024 60000 11144
rect 59200 10480 60000 10600
rect 59200 9936 60000 10056
rect 59200 9392 60000 9512
rect 59200 8848 60000 8968
rect 59200 8304 60000 8424
rect 59200 7760 60000 7880
rect 59200 7216 60000 7336
<< obsm3 >>
rect 4061 72696 59200 78437
rect 4061 72416 59120 72696
rect 4061 72152 59200 72416
rect 4061 71872 59120 72152
rect 4061 71608 59200 71872
rect 4061 71328 59120 71608
rect 4061 71064 59200 71328
rect 4061 70784 59120 71064
rect 4061 70520 59200 70784
rect 4061 70240 59120 70520
rect 4061 69976 59200 70240
rect 4061 69696 59120 69976
rect 4061 69432 59200 69696
rect 4061 69152 59120 69432
rect 4061 68888 59200 69152
rect 4061 68608 59120 68888
rect 4061 68344 59200 68608
rect 4061 68064 59120 68344
rect 4061 67800 59200 68064
rect 4061 67520 59120 67800
rect 4061 67256 59200 67520
rect 4061 66976 59120 67256
rect 4061 66712 59200 66976
rect 4061 66432 59120 66712
rect 4061 66168 59200 66432
rect 4061 65888 59120 66168
rect 4061 65624 59200 65888
rect 4061 65344 59120 65624
rect 4061 65080 59200 65344
rect 4061 64800 59120 65080
rect 4061 64536 59200 64800
rect 4061 64256 59120 64536
rect 4061 63992 59200 64256
rect 4061 63712 59120 63992
rect 4061 63448 59200 63712
rect 4061 63168 59120 63448
rect 4061 62904 59200 63168
rect 4061 62624 59120 62904
rect 4061 62360 59200 62624
rect 4061 62080 59120 62360
rect 4061 61816 59200 62080
rect 4061 61536 59120 61816
rect 4061 61272 59200 61536
rect 4061 60992 59120 61272
rect 4061 60728 59200 60992
rect 4061 60448 59120 60728
rect 4061 60184 59200 60448
rect 4061 59904 59120 60184
rect 4061 59640 59200 59904
rect 4061 59360 59120 59640
rect 4061 59096 59200 59360
rect 4061 58816 59120 59096
rect 4061 58552 59200 58816
rect 4061 58272 59120 58552
rect 4061 58008 59200 58272
rect 4061 57728 59120 58008
rect 4061 57464 59200 57728
rect 4061 57184 59120 57464
rect 4061 56920 59200 57184
rect 4061 56640 59120 56920
rect 4061 56376 59200 56640
rect 4061 56096 59120 56376
rect 4061 55832 59200 56096
rect 4061 55552 59120 55832
rect 4061 55288 59200 55552
rect 4061 55008 59120 55288
rect 4061 54744 59200 55008
rect 4061 54464 59120 54744
rect 4061 54200 59200 54464
rect 4061 53920 59120 54200
rect 4061 53656 59200 53920
rect 4061 53376 59120 53656
rect 4061 53112 59200 53376
rect 4061 52832 59120 53112
rect 4061 52568 59200 52832
rect 4061 52288 59120 52568
rect 4061 52024 59200 52288
rect 4061 51744 59120 52024
rect 4061 51480 59200 51744
rect 4061 51200 59120 51480
rect 4061 50936 59200 51200
rect 4061 50656 59120 50936
rect 4061 50392 59200 50656
rect 4061 50112 59120 50392
rect 4061 49848 59200 50112
rect 4061 49568 59120 49848
rect 4061 49304 59200 49568
rect 4061 49024 59120 49304
rect 4061 48760 59200 49024
rect 4061 48480 59120 48760
rect 4061 48216 59200 48480
rect 4061 47936 59120 48216
rect 4061 47672 59200 47936
rect 4061 47392 59120 47672
rect 4061 47128 59200 47392
rect 4061 46848 59120 47128
rect 4061 46584 59200 46848
rect 4061 46304 59120 46584
rect 4061 46040 59200 46304
rect 4061 45760 59120 46040
rect 4061 45496 59200 45760
rect 4061 45216 59120 45496
rect 4061 44952 59200 45216
rect 4061 44672 59120 44952
rect 4061 44408 59200 44672
rect 4061 44128 59120 44408
rect 4061 43864 59200 44128
rect 4061 43584 59120 43864
rect 4061 43320 59200 43584
rect 4061 43040 59120 43320
rect 4061 42776 59200 43040
rect 4061 42496 59120 42776
rect 4061 42232 59200 42496
rect 4061 41952 59120 42232
rect 4061 41688 59200 41952
rect 4061 41408 59120 41688
rect 4061 41144 59200 41408
rect 4061 40864 59120 41144
rect 4061 40600 59200 40864
rect 4061 40320 59120 40600
rect 4061 40056 59200 40320
rect 4061 39776 59120 40056
rect 4061 39512 59200 39776
rect 4061 39232 59120 39512
rect 4061 38968 59200 39232
rect 4061 38688 59120 38968
rect 4061 38424 59200 38688
rect 4061 38144 59120 38424
rect 4061 37880 59200 38144
rect 4061 37600 59120 37880
rect 4061 37336 59200 37600
rect 4061 37056 59120 37336
rect 4061 36792 59200 37056
rect 4061 36512 59120 36792
rect 4061 36248 59200 36512
rect 4061 35968 59120 36248
rect 4061 35704 59200 35968
rect 4061 35424 59120 35704
rect 4061 35160 59200 35424
rect 4061 34880 59120 35160
rect 4061 34616 59200 34880
rect 4061 34336 59120 34616
rect 4061 34072 59200 34336
rect 4061 33792 59120 34072
rect 4061 33528 59200 33792
rect 4061 33248 59120 33528
rect 4061 32984 59200 33248
rect 4061 32704 59120 32984
rect 4061 32440 59200 32704
rect 4061 32160 59120 32440
rect 4061 31896 59200 32160
rect 4061 31616 59120 31896
rect 4061 31352 59200 31616
rect 4061 31072 59120 31352
rect 4061 30808 59200 31072
rect 4061 30528 59120 30808
rect 4061 30264 59200 30528
rect 4061 29984 59120 30264
rect 4061 29720 59200 29984
rect 4061 29440 59120 29720
rect 4061 29176 59200 29440
rect 4061 28896 59120 29176
rect 4061 28632 59200 28896
rect 4061 28352 59120 28632
rect 4061 28088 59200 28352
rect 4061 27808 59120 28088
rect 4061 27544 59200 27808
rect 4061 27264 59120 27544
rect 4061 27000 59200 27264
rect 4061 26720 59120 27000
rect 4061 26456 59200 26720
rect 4061 26176 59120 26456
rect 4061 25912 59200 26176
rect 4061 25632 59120 25912
rect 4061 25368 59200 25632
rect 4061 25088 59120 25368
rect 4061 24824 59200 25088
rect 4061 24544 59120 24824
rect 4061 24280 59200 24544
rect 4061 24000 59120 24280
rect 4061 23736 59200 24000
rect 4061 23456 59120 23736
rect 4061 23192 59200 23456
rect 4061 22912 59120 23192
rect 4061 22648 59200 22912
rect 4061 22368 59120 22648
rect 4061 22104 59200 22368
rect 4061 21824 59120 22104
rect 4061 21560 59200 21824
rect 4061 21280 59120 21560
rect 4061 21016 59200 21280
rect 4061 20736 59120 21016
rect 4061 20472 59200 20736
rect 4061 20192 59120 20472
rect 4061 19928 59200 20192
rect 4061 19648 59120 19928
rect 4061 19384 59200 19648
rect 4061 19104 59120 19384
rect 4061 18840 59200 19104
rect 4061 18560 59120 18840
rect 4061 18296 59200 18560
rect 4061 18016 59120 18296
rect 4061 17752 59200 18016
rect 4061 17472 59120 17752
rect 4061 17208 59200 17472
rect 4061 16928 59120 17208
rect 4061 16664 59200 16928
rect 4061 16384 59120 16664
rect 4061 16120 59200 16384
rect 4061 15840 59120 16120
rect 4061 15576 59200 15840
rect 4061 15296 59120 15576
rect 4061 15032 59200 15296
rect 4061 14752 59120 15032
rect 4061 14488 59200 14752
rect 4061 14208 59120 14488
rect 4061 13944 59200 14208
rect 4061 13664 59120 13944
rect 4061 13400 59200 13664
rect 4061 13120 59120 13400
rect 4061 12856 59200 13120
rect 4061 12576 59120 12856
rect 4061 12312 59200 12576
rect 4061 12032 59120 12312
rect 4061 11768 59200 12032
rect 4061 11488 59120 11768
rect 4061 11224 59200 11488
rect 4061 10944 59120 11224
rect 4061 10680 59200 10944
rect 4061 10400 59120 10680
rect 4061 10136 59200 10400
rect 4061 9856 59120 10136
rect 4061 9592 59200 9856
rect 4061 9312 59120 9592
rect 4061 9048 59200 9312
rect 4061 8768 59120 9048
rect 4061 8504 59200 8768
rect 4061 8224 59120 8504
rect 4061 7960 59200 8224
rect 4061 7680 59120 7960
rect 4061 7416 59200 7680
rect 4061 7136 59120 7416
rect 4061 2143 59200 7136
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
<< obsm4 >>
rect 8155 77920 38765 78437
rect 8155 2483 19488 77920
rect 19968 2483 34848 77920
rect 35328 2483 38765 77920
<< labels >>
rlabel metal2 s 1398 0 1454 800 6 inner_clock
port 1 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 inner_disable
port 2 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 inner_embed_mode
port 3 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 inner_ext_irq
port 4 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 inner_reset
port 5 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 inner_wb_4_burst
port 6 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 inner_wb_8_burst
port 7 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 inner_wb_ack
port 8 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 inner_wb_adr[0]
port 9 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 inner_wb_adr[10]
port 10 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 inner_wb_adr[11]
port 11 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 inner_wb_adr[12]
port 12 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 inner_wb_adr[13]
port 13 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 inner_wb_adr[14]
port 14 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 inner_wb_adr[15]
port 15 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 inner_wb_adr[16]
port 16 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 inner_wb_adr[17]
port 17 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 inner_wb_adr[18]
port 18 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 inner_wb_adr[19]
port 19 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 inner_wb_adr[1]
port 20 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 inner_wb_adr[20]
port 21 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 inner_wb_adr[21]
port 22 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 inner_wb_adr[22]
port 23 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 inner_wb_adr[23]
port 24 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 inner_wb_adr[2]
port 25 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 inner_wb_adr[3]
port 26 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 inner_wb_adr[4]
port 27 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 inner_wb_adr[5]
port 28 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 inner_wb_adr[6]
port 29 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 inner_wb_adr[7]
port 30 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 inner_wb_adr[8]
port 31 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 inner_wb_adr[9]
port 32 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 inner_wb_cyc
port 33 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 inner_wb_err
port 34 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 inner_wb_i_dat[0]
port 35 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 inner_wb_i_dat[10]
port 36 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 inner_wb_i_dat[11]
port 37 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 inner_wb_i_dat[12]
port 38 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 inner_wb_i_dat[13]
port 39 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 inner_wb_i_dat[14]
port 40 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 inner_wb_i_dat[15]
port 41 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 inner_wb_i_dat[1]
port 42 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 inner_wb_i_dat[2]
port 43 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 inner_wb_i_dat[3]
port 44 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 inner_wb_i_dat[4]
port 45 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 inner_wb_i_dat[5]
port 46 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 inner_wb_i_dat[6]
port 47 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 inner_wb_i_dat[7]
port 48 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 inner_wb_i_dat[8]
port 49 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 inner_wb_i_dat[9]
port 50 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 inner_wb_o_dat[0]
port 51 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 inner_wb_o_dat[10]
port 52 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 inner_wb_o_dat[11]
port 53 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 inner_wb_o_dat[12]
port 54 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 inner_wb_o_dat[13]
port 55 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 inner_wb_o_dat[14]
port 56 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 inner_wb_o_dat[15]
port 57 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 inner_wb_o_dat[1]
port 58 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 inner_wb_o_dat[2]
port 59 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 inner_wb_o_dat[3]
port 60 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 inner_wb_o_dat[4]
port 61 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 inner_wb_o_dat[5]
port 62 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 inner_wb_o_dat[6]
port 63 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 inner_wb_o_dat[7]
port 64 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 inner_wb_o_dat[8]
port 65 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 inner_wb_o_dat[9]
port 66 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 inner_wb_sel[0]
port 67 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 inner_wb_sel[1]
port 68 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 inner_wb_stb
port 69 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 inner_wb_we
port 70 nsew signal input
rlabel metal3 s 59200 9936 60000 10056 6 iram1_addr[0]
port 71 nsew signal output
rlabel metal3 s 59200 13200 60000 13320 6 iram1_addr[1]
port 72 nsew signal output
rlabel metal3 s 59200 16464 60000 16584 6 iram1_addr[2]
port 73 nsew signal output
rlabel metal3 s 59200 19728 60000 19848 6 iram1_addr[3]
port 74 nsew signal output
rlabel metal3 s 59200 22992 60000 23112 6 iram1_addr[4]
port 75 nsew signal output
rlabel metal3 s 59200 25712 60000 25832 6 iram1_addr[5]
port 76 nsew signal output
rlabel metal3 s 59200 28432 60000 28552 6 iram1_addr[6]
port 77 nsew signal output
rlabel metal3 s 59200 31152 60000 31272 6 iram1_addr[7]
port 78 nsew signal output
rlabel metal3 s 59200 7216 60000 7336 6 iram1_clk
port 79 nsew signal input
rlabel metal3 s 59200 7760 60000 7880 6 iram1_csb
port 80 nsew signal input
rlabel metal3 s 59200 10480 60000 10600 6 iram1_dout[0]
port 81 nsew signal input
rlabel metal3 s 59200 37136 60000 37256 6 iram1_dout[10]
port 82 nsew signal input
rlabel metal3 s 59200 38768 60000 38888 6 iram1_dout[11]
port 83 nsew signal input
rlabel metal3 s 59200 40400 60000 40520 6 iram1_dout[12]
port 84 nsew signal input
rlabel metal3 s 59200 42032 60000 42152 6 iram1_dout[13]
port 85 nsew signal input
rlabel metal3 s 59200 43664 60000 43784 6 iram1_dout[14]
port 86 nsew signal input
rlabel metal3 s 59200 45296 60000 45416 6 iram1_dout[15]
port 87 nsew signal input
rlabel metal3 s 59200 46928 60000 47048 6 iram1_dout[16]
port 88 nsew signal input
rlabel metal3 s 59200 48560 60000 48680 6 iram1_dout[17]
port 89 nsew signal input
rlabel metal3 s 59200 50192 60000 50312 6 iram1_dout[18]
port 90 nsew signal input
rlabel metal3 s 59200 51824 60000 51944 6 iram1_dout[19]
port 91 nsew signal input
rlabel metal3 s 59200 13744 60000 13864 6 iram1_dout[1]
port 92 nsew signal input
rlabel metal3 s 59200 53456 60000 53576 6 iram1_dout[20]
port 93 nsew signal input
rlabel metal3 s 59200 55088 60000 55208 6 iram1_dout[21]
port 94 nsew signal input
rlabel metal3 s 59200 56720 60000 56840 6 iram1_dout[22]
port 95 nsew signal input
rlabel metal3 s 59200 58352 60000 58472 6 iram1_dout[23]
port 96 nsew signal input
rlabel metal3 s 59200 59984 60000 60104 6 iram1_dout[24]
port 97 nsew signal input
rlabel metal3 s 59200 61616 60000 61736 6 iram1_dout[25]
port 98 nsew signal input
rlabel metal3 s 59200 63248 60000 63368 6 iram1_dout[26]
port 99 nsew signal input
rlabel metal3 s 59200 64880 60000 65000 6 iram1_dout[27]
port 100 nsew signal input
rlabel metal3 s 59200 66512 60000 66632 6 iram1_dout[28]
port 101 nsew signal input
rlabel metal3 s 59200 68144 60000 68264 6 iram1_dout[29]
port 102 nsew signal input
rlabel metal3 s 59200 17008 60000 17128 6 iram1_dout[2]
port 103 nsew signal input
rlabel metal3 s 59200 69776 60000 69896 6 iram1_dout[30]
port 104 nsew signal input
rlabel metal3 s 59200 71408 60000 71528 6 iram1_dout[31]
port 105 nsew signal input
rlabel metal3 s 59200 20272 60000 20392 6 iram1_dout[3]
port 106 nsew signal input
rlabel metal3 s 59200 23536 60000 23656 6 iram1_dout[4]
port 107 nsew signal input
rlabel metal3 s 59200 26256 60000 26376 6 iram1_dout[5]
port 108 nsew signal input
rlabel metal3 s 59200 28976 60000 29096 6 iram1_dout[6]
port 109 nsew signal input
rlabel metal3 s 59200 31696 60000 31816 6 iram1_dout[7]
port 110 nsew signal input
rlabel metal3 s 59200 33872 60000 33992 6 iram1_dout[8]
port 111 nsew signal input
rlabel metal3 s 59200 35504 60000 35624 6 iram1_dout[9]
port 112 nsew signal input
rlabel metal3 s 59200 11024 60000 11144 6 iram_addr[0]
port 113 nsew signal output
rlabel metal3 s 59200 14288 60000 14408 6 iram_addr[1]
port 114 nsew signal output
rlabel metal3 s 59200 17552 60000 17672 6 iram_addr[2]
port 115 nsew signal output
rlabel metal3 s 59200 20816 60000 20936 6 iram_addr[3]
port 116 nsew signal output
rlabel metal3 s 59200 24080 60000 24200 6 iram_addr[4]
port 117 nsew signal output
rlabel metal3 s 59200 26800 60000 26920 6 iram_addr[5]
port 118 nsew signal output
rlabel metal3 s 59200 29520 60000 29640 6 iram_addr[6]
port 119 nsew signal output
rlabel metal3 s 59200 32240 60000 32360 6 iram_addr[7]
port 120 nsew signal output
rlabel metal3 s 59200 8304 60000 8424 6 iram_clk
port 121 nsew signal output
rlabel metal3 s 59200 8848 60000 8968 6 iram_csb
port 122 nsew signal output
rlabel metal3 s 59200 11568 60000 11688 6 iram_i_data[0]
port 123 nsew signal output
rlabel metal3 s 59200 37680 60000 37800 6 iram_i_data[10]
port 124 nsew signal output
rlabel metal3 s 59200 39312 60000 39432 6 iram_i_data[11]
port 125 nsew signal output
rlabel metal3 s 59200 40944 60000 41064 6 iram_i_data[12]
port 126 nsew signal output
rlabel metal3 s 59200 42576 60000 42696 6 iram_i_data[13]
port 127 nsew signal output
rlabel metal3 s 59200 44208 60000 44328 6 iram_i_data[14]
port 128 nsew signal output
rlabel metal3 s 59200 45840 60000 45960 6 iram_i_data[15]
port 129 nsew signal output
rlabel metal3 s 59200 47472 60000 47592 6 iram_i_data[16]
port 130 nsew signal output
rlabel metal3 s 59200 49104 60000 49224 6 iram_i_data[17]
port 131 nsew signal output
rlabel metal3 s 59200 50736 60000 50856 6 iram_i_data[18]
port 132 nsew signal output
rlabel metal3 s 59200 52368 60000 52488 6 iram_i_data[19]
port 133 nsew signal output
rlabel metal3 s 59200 14832 60000 14952 6 iram_i_data[1]
port 134 nsew signal output
rlabel metal3 s 59200 54000 60000 54120 6 iram_i_data[20]
port 135 nsew signal output
rlabel metal3 s 59200 55632 60000 55752 6 iram_i_data[21]
port 136 nsew signal output
rlabel metal3 s 59200 57264 60000 57384 6 iram_i_data[22]
port 137 nsew signal output
rlabel metal3 s 59200 58896 60000 59016 6 iram_i_data[23]
port 138 nsew signal output
rlabel metal3 s 59200 60528 60000 60648 6 iram_i_data[24]
port 139 nsew signal output
rlabel metal3 s 59200 62160 60000 62280 6 iram_i_data[25]
port 140 nsew signal output
rlabel metal3 s 59200 63792 60000 63912 6 iram_i_data[26]
port 141 nsew signal output
rlabel metal3 s 59200 65424 60000 65544 6 iram_i_data[27]
port 142 nsew signal output
rlabel metal3 s 59200 67056 60000 67176 6 iram_i_data[28]
port 143 nsew signal output
rlabel metal3 s 59200 68688 60000 68808 6 iram_i_data[29]
port 144 nsew signal output
rlabel metal3 s 59200 18096 60000 18216 6 iram_i_data[2]
port 145 nsew signal output
rlabel metal3 s 59200 70320 60000 70440 6 iram_i_data[30]
port 146 nsew signal output
rlabel metal3 s 59200 71952 60000 72072 6 iram_i_data[31]
port 147 nsew signal output
rlabel metal3 s 59200 21360 60000 21480 6 iram_i_data[3]
port 148 nsew signal output
rlabel metal3 s 59200 24624 60000 24744 6 iram_i_data[4]
port 149 nsew signal output
rlabel metal3 s 59200 27344 60000 27464 6 iram_i_data[5]
port 150 nsew signal output
rlabel metal3 s 59200 30064 60000 30184 6 iram_i_data[6]
port 151 nsew signal output
rlabel metal3 s 59200 32784 60000 32904 6 iram_i_data[7]
port 152 nsew signal output
rlabel metal3 s 59200 34416 60000 34536 6 iram_i_data[8]
port 153 nsew signal output
rlabel metal3 s 59200 36048 60000 36168 6 iram_i_data[9]
port 154 nsew signal output
rlabel metal3 s 59200 12112 60000 12232 6 iram_o_data[0]
port 155 nsew signal input
rlabel metal3 s 59200 38224 60000 38344 6 iram_o_data[10]
port 156 nsew signal input
rlabel metal3 s 59200 39856 60000 39976 6 iram_o_data[11]
port 157 nsew signal input
rlabel metal3 s 59200 41488 60000 41608 6 iram_o_data[12]
port 158 nsew signal input
rlabel metal3 s 59200 43120 60000 43240 6 iram_o_data[13]
port 159 nsew signal input
rlabel metal3 s 59200 44752 60000 44872 6 iram_o_data[14]
port 160 nsew signal input
rlabel metal3 s 59200 46384 60000 46504 6 iram_o_data[15]
port 161 nsew signal input
rlabel metal3 s 59200 48016 60000 48136 6 iram_o_data[16]
port 162 nsew signal input
rlabel metal3 s 59200 49648 60000 49768 6 iram_o_data[17]
port 163 nsew signal input
rlabel metal3 s 59200 51280 60000 51400 6 iram_o_data[18]
port 164 nsew signal input
rlabel metal3 s 59200 52912 60000 53032 6 iram_o_data[19]
port 165 nsew signal input
rlabel metal3 s 59200 15376 60000 15496 6 iram_o_data[1]
port 166 nsew signal input
rlabel metal3 s 59200 54544 60000 54664 6 iram_o_data[20]
port 167 nsew signal input
rlabel metal3 s 59200 56176 60000 56296 6 iram_o_data[21]
port 168 nsew signal input
rlabel metal3 s 59200 57808 60000 57928 6 iram_o_data[22]
port 169 nsew signal input
rlabel metal3 s 59200 59440 60000 59560 6 iram_o_data[23]
port 170 nsew signal input
rlabel metal3 s 59200 61072 60000 61192 6 iram_o_data[24]
port 171 nsew signal input
rlabel metal3 s 59200 62704 60000 62824 6 iram_o_data[25]
port 172 nsew signal input
rlabel metal3 s 59200 64336 60000 64456 6 iram_o_data[26]
port 173 nsew signal input
rlabel metal3 s 59200 65968 60000 66088 6 iram_o_data[27]
port 174 nsew signal input
rlabel metal3 s 59200 67600 60000 67720 6 iram_o_data[28]
port 175 nsew signal input
rlabel metal3 s 59200 69232 60000 69352 6 iram_o_data[29]
port 176 nsew signal input
rlabel metal3 s 59200 18640 60000 18760 6 iram_o_data[2]
port 177 nsew signal input
rlabel metal3 s 59200 70864 60000 70984 6 iram_o_data[30]
port 178 nsew signal input
rlabel metal3 s 59200 72496 60000 72616 6 iram_o_data[31]
port 179 nsew signal input
rlabel metal3 s 59200 21904 60000 22024 6 iram_o_data[3]
port 180 nsew signal input
rlabel metal3 s 59200 25168 60000 25288 6 iram_o_data[4]
port 181 nsew signal input
rlabel metal3 s 59200 27888 60000 28008 6 iram_o_data[5]
port 182 nsew signal input
rlabel metal3 s 59200 30608 60000 30728 6 iram_o_data[6]
port 183 nsew signal input
rlabel metal3 s 59200 33328 60000 33448 6 iram_o_data[7]
port 184 nsew signal input
rlabel metal3 s 59200 34960 60000 35080 6 iram_o_data[8]
port 185 nsew signal input
rlabel metal3 s 59200 36592 60000 36712 6 iram_o_data[9]
port 186 nsew signal input
rlabel metal3 s 59200 12656 60000 12776 6 iram_w_mask[0]
port 187 nsew signal output
rlabel metal3 s 59200 15920 60000 16040 6 iram_w_mask[1]
port 188 nsew signal output
rlabel metal3 s 59200 19184 60000 19304 6 iram_w_mask[2]
port 189 nsew signal output
rlabel metal3 s 59200 22448 60000 22568 6 iram_w_mask[3]
port 190 nsew signal output
rlabel metal3 s 59200 9392 60000 9512 6 iram_we
port 191 nsew signal output
rlabel metal2 s 57610 79200 57666 80000 6 irq[0]
port 192 nsew signal output
rlabel metal2 s 57702 79200 57758 80000 6 irq[1]
port 193 nsew signal output
rlabel metal2 s 57794 79200 57850 80000 6 irq[2]
port 194 nsew signal output
rlabel metal2 s 22282 79200 22338 80000 6 la_data_in[0]
port 195 nsew signal input
rlabel metal2 s 49882 79200 49938 80000 6 la_data_in[100]
port 196 nsew signal input
rlabel metal2 s 50158 79200 50214 80000 6 la_data_in[101]
port 197 nsew signal input
rlabel metal2 s 50434 79200 50490 80000 6 la_data_in[102]
port 198 nsew signal input
rlabel metal2 s 50710 79200 50766 80000 6 la_data_in[103]
port 199 nsew signal input
rlabel metal2 s 50986 79200 51042 80000 6 la_data_in[104]
port 200 nsew signal input
rlabel metal2 s 51262 79200 51318 80000 6 la_data_in[105]
port 201 nsew signal input
rlabel metal2 s 51538 79200 51594 80000 6 la_data_in[106]
port 202 nsew signal input
rlabel metal2 s 51814 79200 51870 80000 6 la_data_in[107]
port 203 nsew signal input
rlabel metal2 s 52090 79200 52146 80000 6 la_data_in[108]
port 204 nsew signal input
rlabel metal2 s 52366 79200 52422 80000 6 la_data_in[109]
port 205 nsew signal input
rlabel metal2 s 25042 79200 25098 80000 6 la_data_in[10]
port 206 nsew signal input
rlabel metal2 s 52642 79200 52698 80000 6 la_data_in[110]
port 207 nsew signal input
rlabel metal2 s 52918 79200 52974 80000 6 la_data_in[111]
port 208 nsew signal input
rlabel metal2 s 53194 79200 53250 80000 6 la_data_in[112]
port 209 nsew signal input
rlabel metal2 s 53470 79200 53526 80000 6 la_data_in[113]
port 210 nsew signal input
rlabel metal2 s 53746 79200 53802 80000 6 la_data_in[114]
port 211 nsew signal input
rlabel metal2 s 54022 79200 54078 80000 6 la_data_in[115]
port 212 nsew signal input
rlabel metal2 s 54298 79200 54354 80000 6 la_data_in[116]
port 213 nsew signal input
rlabel metal2 s 54574 79200 54630 80000 6 la_data_in[117]
port 214 nsew signal input
rlabel metal2 s 54850 79200 54906 80000 6 la_data_in[118]
port 215 nsew signal input
rlabel metal2 s 55126 79200 55182 80000 6 la_data_in[119]
port 216 nsew signal input
rlabel metal2 s 25318 79200 25374 80000 6 la_data_in[11]
port 217 nsew signal input
rlabel metal2 s 55402 79200 55458 80000 6 la_data_in[120]
port 218 nsew signal input
rlabel metal2 s 55678 79200 55734 80000 6 la_data_in[121]
port 219 nsew signal input
rlabel metal2 s 55954 79200 56010 80000 6 la_data_in[122]
port 220 nsew signal input
rlabel metal2 s 56230 79200 56286 80000 6 la_data_in[123]
port 221 nsew signal input
rlabel metal2 s 56506 79200 56562 80000 6 la_data_in[124]
port 222 nsew signal input
rlabel metal2 s 56782 79200 56838 80000 6 la_data_in[125]
port 223 nsew signal input
rlabel metal2 s 57058 79200 57114 80000 6 la_data_in[126]
port 224 nsew signal input
rlabel metal2 s 57334 79200 57390 80000 6 la_data_in[127]
port 225 nsew signal input
rlabel metal2 s 25594 79200 25650 80000 6 la_data_in[12]
port 226 nsew signal input
rlabel metal2 s 25870 79200 25926 80000 6 la_data_in[13]
port 227 nsew signal input
rlabel metal2 s 26146 79200 26202 80000 6 la_data_in[14]
port 228 nsew signal input
rlabel metal2 s 26422 79200 26478 80000 6 la_data_in[15]
port 229 nsew signal input
rlabel metal2 s 26698 79200 26754 80000 6 la_data_in[16]
port 230 nsew signal input
rlabel metal2 s 26974 79200 27030 80000 6 la_data_in[17]
port 231 nsew signal input
rlabel metal2 s 27250 79200 27306 80000 6 la_data_in[18]
port 232 nsew signal input
rlabel metal2 s 27526 79200 27582 80000 6 la_data_in[19]
port 233 nsew signal input
rlabel metal2 s 22558 79200 22614 80000 6 la_data_in[1]
port 234 nsew signal input
rlabel metal2 s 27802 79200 27858 80000 6 la_data_in[20]
port 235 nsew signal input
rlabel metal2 s 28078 79200 28134 80000 6 la_data_in[21]
port 236 nsew signal input
rlabel metal2 s 28354 79200 28410 80000 6 la_data_in[22]
port 237 nsew signal input
rlabel metal2 s 28630 79200 28686 80000 6 la_data_in[23]
port 238 nsew signal input
rlabel metal2 s 28906 79200 28962 80000 6 la_data_in[24]
port 239 nsew signal input
rlabel metal2 s 29182 79200 29238 80000 6 la_data_in[25]
port 240 nsew signal input
rlabel metal2 s 29458 79200 29514 80000 6 la_data_in[26]
port 241 nsew signal input
rlabel metal2 s 29734 79200 29790 80000 6 la_data_in[27]
port 242 nsew signal input
rlabel metal2 s 30010 79200 30066 80000 6 la_data_in[28]
port 243 nsew signal input
rlabel metal2 s 30286 79200 30342 80000 6 la_data_in[29]
port 244 nsew signal input
rlabel metal2 s 22834 79200 22890 80000 6 la_data_in[2]
port 245 nsew signal input
rlabel metal2 s 30562 79200 30618 80000 6 la_data_in[30]
port 246 nsew signal input
rlabel metal2 s 30838 79200 30894 80000 6 la_data_in[31]
port 247 nsew signal input
rlabel metal2 s 31114 79200 31170 80000 6 la_data_in[32]
port 248 nsew signal input
rlabel metal2 s 31390 79200 31446 80000 6 la_data_in[33]
port 249 nsew signal input
rlabel metal2 s 31666 79200 31722 80000 6 la_data_in[34]
port 250 nsew signal input
rlabel metal2 s 31942 79200 31998 80000 6 la_data_in[35]
port 251 nsew signal input
rlabel metal2 s 32218 79200 32274 80000 6 la_data_in[36]
port 252 nsew signal input
rlabel metal2 s 32494 79200 32550 80000 6 la_data_in[37]
port 253 nsew signal input
rlabel metal2 s 32770 79200 32826 80000 6 la_data_in[38]
port 254 nsew signal input
rlabel metal2 s 33046 79200 33102 80000 6 la_data_in[39]
port 255 nsew signal input
rlabel metal2 s 23110 79200 23166 80000 6 la_data_in[3]
port 256 nsew signal input
rlabel metal2 s 33322 79200 33378 80000 6 la_data_in[40]
port 257 nsew signal input
rlabel metal2 s 33598 79200 33654 80000 6 la_data_in[41]
port 258 nsew signal input
rlabel metal2 s 33874 79200 33930 80000 6 la_data_in[42]
port 259 nsew signal input
rlabel metal2 s 34150 79200 34206 80000 6 la_data_in[43]
port 260 nsew signal input
rlabel metal2 s 34426 79200 34482 80000 6 la_data_in[44]
port 261 nsew signal input
rlabel metal2 s 34702 79200 34758 80000 6 la_data_in[45]
port 262 nsew signal input
rlabel metal2 s 34978 79200 35034 80000 6 la_data_in[46]
port 263 nsew signal input
rlabel metal2 s 35254 79200 35310 80000 6 la_data_in[47]
port 264 nsew signal input
rlabel metal2 s 35530 79200 35586 80000 6 la_data_in[48]
port 265 nsew signal input
rlabel metal2 s 35806 79200 35862 80000 6 la_data_in[49]
port 266 nsew signal input
rlabel metal2 s 23386 79200 23442 80000 6 la_data_in[4]
port 267 nsew signal input
rlabel metal2 s 36082 79200 36138 80000 6 la_data_in[50]
port 268 nsew signal input
rlabel metal2 s 36358 79200 36414 80000 6 la_data_in[51]
port 269 nsew signal input
rlabel metal2 s 36634 79200 36690 80000 6 la_data_in[52]
port 270 nsew signal input
rlabel metal2 s 36910 79200 36966 80000 6 la_data_in[53]
port 271 nsew signal input
rlabel metal2 s 37186 79200 37242 80000 6 la_data_in[54]
port 272 nsew signal input
rlabel metal2 s 37462 79200 37518 80000 6 la_data_in[55]
port 273 nsew signal input
rlabel metal2 s 37738 79200 37794 80000 6 la_data_in[56]
port 274 nsew signal input
rlabel metal2 s 38014 79200 38070 80000 6 la_data_in[57]
port 275 nsew signal input
rlabel metal2 s 38290 79200 38346 80000 6 la_data_in[58]
port 276 nsew signal input
rlabel metal2 s 38566 79200 38622 80000 6 la_data_in[59]
port 277 nsew signal input
rlabel metal2 s 23662 79200 23718 80000 6 la_data_in[5]
port 278 nsew signal input
rlabel metal2 s 38842 79200 38898 80000 6 la_data_in[60]
port 279 nsew signal input
rlabel metal2 s 39118 79200 39174 80000 6 la_data_in[61]
port 280 nsew signal input
rlabel metal2 s 39394 79200 39450 80000 6 la_data_in[62]
port 281 nsew signal input
rlabel metal2 s 39670 79200 39726 80000 6 la_data_in[63]
port 282 nsew signal input
rlabel metal2 s 39946 79200 40002 80000 6 la_data_in[64]
port 283 nsew signal input
rlabel metal2 s 40222 79200 40278 80000 6 la_data_in[65]
port 284 nsew signal input
rlabel metal2 s 40498 79200 40554 80000 6 la_data_in[66]
port 285 nsew signal input
rlabel metal2 s 40774 79200 40830 80000 6 la_data_in[67]
port 286 nsew signal input
rlabel metal2 s 41050 79200 41106 80000 6 la_data_in[68]
port 287 nsew signal input
rlabel metal2 s 41326 79200 41382 80000 6 la_data_in[69]
port 288 nsew signal input
rlabel metal2 s 23938 79200 23994 80000 6 la_data_in[6]
port 289 nsew signal input
rlabel metal2 s 41602 79200 41658 80000 6 la_data_in[70]
port 290 nsew signal input
rlabel metal2 s 41878 79200 41934 80000 6 la_data_in[71]
port 291 nsew signal input
rlabel metal2 s 42154 79200 42210 80000 6 la_data_in[72]
port 292 nsew signal input
rlabel metal2 s 42430 79200 42486 80000 6 la_data_in[73]
port 293 nsew signal input
rlabel metal2 s 42706 79200 42762 80000 6 la_data_in[74]
port 294 nsew signal input
rlabel metal2 s 42982 79200 43038 80000 6 la_data_in[75]
port 295 nsew signal input
rlabel metal2 s 43258 79200 43314 80000 6 la_data_in[76]
port 296 nsew signal input
rlabel metal2 s 43534 79200 43590 80000 6 la_data_in[77]
port 297 nsew signal input
rlabel metal2 s 43810 79200 43866 80000 6 la_data_in[78]
port 298 nsew signal input
rlabel metal2 s 44086 79200 44142 80000 6 la_data_in[79]
port 299 nsew signal input
rlabel metal2 s 24214 79200 24270 80000 6 la_data_in[7]
port 300 nsew signal input
rlabel metal2 s 44362 79200 44418 80000 6 la_data_in[80]
port 301 nsew signal input
rlabel metal2 s 44638 79200 44694 80000 6 la_data_in[81]
port 302 nsew signal input
rlabel metal2 s 44914 79200 44970 80000 6 la_data_in[82]
port 303 nsew signal input
rlabel metal2 s 45190 79200 45246 80000 6 la_data_in[83]
port 304 nsew signal input
rlabel metal2 s 45466 79200 45522 80000 6 la_data_in[84]
port 305 nsew signal input
rlabel metal2 s 45742 79200 45798 80000 6 la_data_in[85]
port 306 nsew signal input
rlabel metal2 s 46018 79200 46074 80000 6 la_data_in[86]
port 307 nsew signal input
rlabel metal2 s 46294 79200 46350 80000 6 la_data_in[87]
port 308 nsew signal input
rlabel metal2 s 46570 79200 46626 80000 6 la_data_in[88]
port 309 nsew signal input
rlabel metal2 s 46846 79200 46902 80000 6 la_data_in[89]
port 310 nsew signal input
rlabel metal2 s 24490 79200 24546 80000 6 la_data_in[8]
port 311 nsew signal input
rlabel metal2 s 47122 79200 47178 80000 6 la_data_in[90]
port 312 nsew signal input
rlabel metal2 s 47398 79200 47454 80000 6 la_data_in[91]
port 313 nsew signal input
rlabel metal2 s 47674 79200 47730 80000 6 la_data_in[92]
port 314 nsew signal input
rlabel metal2 s 47950 79200 48006 80000 6 la_data_in[93]
port 315 nsew signal input
rlabel metal2 s 48226 79200 48282 80000 6 la_data_in[94]
port 316 nsew signal input
rlabel metal2 s 48502 79200 48558 80000 6 la_data_in[95]
port 317 nsew signal input
rlabel metal2 s 48778 79200 48834 80000 6 la_data_in[96]
port 318 nsew signal input
rlabel metal2 s 49054 79200 49110 80000 6 la_data_in[97]
port 319 nsew signal input
rlabel metal2 s 49330 79200 49386 80000 6 la_data_in[98]
port 320 nsew signal input
rlabel metal2 s 49606 79200 49662 80000 6 la_data_in[99]
port 321 nsew signal input
rlabel metal2 s 24766 79200 24822 80000 6 la_data_in[9]
port 322 nsew signal input
rlabel metal2 s 22374 79200 22430 80000 6 la_data_out[0]
port 323 nsew signal output
rlabel metal2 s 49974 79200 50030 80000 6 la_data_out[100]
port 324 nsew signal output
rlabel metal2 s 50250 79200 50306 80000 6 la_data_out[101]
port 325 nsew signal output
rlabel metal2 s 50526 79200 50582 80000 6 la_data_out[102]
port 326 nsew signal output
rlabel metal2 s 50802 79200 50858 80000 6 la_data_out[103]
port 327 nsew signal output
rlabel metal2 s 51078 79200 51134 80000 6 la_data_out[104]
port 328 nsew signal output
rlabel metal2 s 51354 79200 51410 80000 6 la_data_out[105]
port 329 nsew signal output
rlabel metal2 s 51630 79200 51686 80000 6 la_data_out[106]
port 330 nsew signal output
rlabel metal2 s 51906 79200 51962 80000 6 la_data_out[107]
port 331 nsew signal output
rlabel metal2 s 52182 79200 52238 80000 6 la_data_out[108]
port 332 nsew signal output
rlabel metal2 s 52458 79200 52514 80000 6 la_data_out[109]
port 333 nsew signal output
rlabel metal2 s 25134 79200 25190 80000 6 la_data_out[10]
port 334 nsew signal output
rlabel metal2 s 52734 79200 52790 80000 6 la_data_out[110]
port 335 nsew signal output
rlabel metal2 s 53010 79200 53066 80000 6 la_data_out[111]
port 336 nsew signal output
rlabel metal2 s 53286 79200 53342 80000 6 la_data_out[112]
port 337 nsew signal output
rlabel metal2 s 53562 79200 53618 80000 6 la_data_out[113]
port 338 nsew signal output
rlabel metal2 s 53838 79200 53894 80000 6 la_data_out[114]
port 339 nsew signal output
rlabel metal2 s 54114 79200 54170 80000 6 la_data_out[115]
port 340 nsew signal output
rlabel metal2 s 54390 79200 54446 80000 6 la_data_out[116]
port 341 nsew signal output
rlabel metal2 s 54666 79200 54722 80000 6 la_data_out[117]
port 342 nsew signal output
rlabel metal2 s 54942 79200 54998 80000 6 la_data_out[118]
port 343 nsew signal output
rlabel metal2 s 55218 79200 55274 80000 6 la_data_out[119]
port 344 nsew signal output
rlabel metal2 s 25410 79200 25466 80000 6 la_data_out[11]
port 345 nsew signal output
rlabel metal2 s 55494 79200 55550 80000 6 la_data_out[120]
port 346 nsew signal output
rlabel metal2 s 55770 79200 55826 80000 6 la_data_out[121]
port 347 nsew signal output
rlabel metal2 s 56046 79200 56102 80000 6 la_data_out[122]
port 348 nsew signal output
rlabel metal2 s 56322 79200 56378 80000 6 la_data_out[123]
port 349 nsew signal output
rlabel metal2 s 56598 79200 56654 80000 6 la_data_out[124]
port 350 nsew signal output
rlabel metal2 s 56874 79200 56930 80000 6 la_data_out[125]
port 351 nsew signal output
rlabel metal2 s 57150 79200 57206 80000 6 la_data_out[126]
port 352 nsew signal output
rlabel metal2 s 57426 79200 57482 80000 6 la_data_out[127]
port 353 nsew signal output
rlabel metal2 s 25686 79200 25742 80000 6 la_data_out[12]
port 354 nsew signal output
rlabel metal2 s 25962 79200 26018 80000 6 la_data_out[13]
port 355 nsew signal output
rlabel metal2 s 26238 79200 26294 80000 6 la_data_out[14]
port 356 nsew signal output
rlabel metal2 s 26514 79200 26570 80000 6 la_data_out[15]
port 357 nsew signal output
rlabel metal2 s 26790 79200 26846 80000 6 la_data_out[16]
port 358 nsew signal output
rlabel metal2 s 27066 79200 27122 80000 6 la_data_out[17]
port 359 nsew signal output
rlabel metal2 s 27342 79200 27398 80000 6 la_data_out[18]
port 360 nsew signal output
rlabel metal2 s 27618 79200 27674 80000 6 la_data_out[19]
port 361 nsew signal output
rlabel metal2 s 22650 79200 22706 80000 6 la_data_out[1]
port 362 nsew signal output
rlabel metal2 s 27894 79200 27950 80000 6 la_data_out[20]
port 363 nsew signal output
rlabel metal2 s 28170 79200 28226 80000 6 la_data_out[21]
port 364 nsew signal output
rlabel metal2 s 28446 79200 28502 80000 6 la_data_out[22]
port 365 nsew signal output
rlabel metal2 s 28722 79200 28778 80000 6 la_data_out[23]
port 366 nsew signal output
rlabel metal2 s 28998 79200 29054 80000 6 la_data_out[24]
port 367 nsew signal output
rlabel metal2 s 29274 79200 29330 80000 6 la_data_out[25]
port 368 nsew signal output
rlabel metal2 s 29550 79200 29606 80000 6 la_data_out[26]
port 369 nsew signal output
rlabel metal2 s 29826 79200 29882 80000 6 la_data_out[27]
port 370 nsew signal output
rlabel metal2 s 30102 79200 30158 80000 6 la_data_out[28]
port 371 nsew signal output
rlabel metal2 s 30378 79200 30434 80000 6 la_data_out[29]
port 372 nsew signal output
rlabel metal2 s 22926 79200 22982 80000 6 la_data_out[2]
port 373 nsew signal output
rlabel metal2 s 30654 79200 30710 80000 6 la_data_out[30]
port 374 nsew signal output
rlabel metal2 s 30930 79200 30986 80000 6 la_data_out[31]
port 375 nsew signal output
rlabel metal2 s 31206 79200 31262 80000 6 la_data_out[32]
port 376 nsew signal output
rlabel metal2 s 31482 79200 31538 80000 6 la_data_out[33]
port 377 nsew signal output
rlabel metal2 s 31758 79200 31814 80000 6 la_data_out[34]
port 378 nsew signal output
rlabel metal2 s 32034 79200 32090 80000 6 la_data_out[35]
port 379 nsew signal output
rlabel metal2 s 32310 79200 32366 80000 6 la_data_out[36]
port 380 nsew signal output
rlabel metal2 s 32586 79200 32642 80000 6 la_data_out[37]
port 381 nsew signal output
rlabel metal2 s 32862 79200 32918 80000 6 la_data_out[38]
port 382 nsew signal output
rlabel metal2 s 33138 79200 33194 80000 6 la_data_out[39]
port 383 nsew signal output
rlabel metal2 s 23202 79200 23258 80000 6 la_data_out[3]
port 384 nsew signal output
rlabel metal2 s 33414 79200 33470 80000 6 la_data_out[40]
port 385 nsew signal output
rlabel metal2 s 33690 79200 33746 80000 6 la_data_out[41]
port 386 nsew signal output
rlabel metal2 s 33966 79200 34022 80000 6 la_data_out[42]
port 387 nsew signal output
rlabel metal2 s 34242 79200 34298 80000 6 la_data_out[43]
port 388 nsew signal output
rlabel metal2 s 34518 79200 34574 80000 6 la_data_out[44]
port 389 nsew signal output
rlabel metal2 s 34794 79200 34850 80000 6 la_data_out[45]
port 390 nsew signal output
rlabel metal2 s 35070 79200 35126 80000 6 la_data_out[46]
port 391 nsew signal output
rlabel metal2 s 35346 79200 35402 80000 6 la_data_out[47]
port 392 nsew signal output
rlabel metal2 s 35622 79200 35678 80000 6 la_data_out[48]
port 393 nsew signal output
rlabel metal2 s 35898 79200 35954 80000 6 la_data_out[49]
port 394 nsew signal output
rlabel metal2 s 23478 79200 23534 80000 6 la_data_out[4]
port 395 nsew signal output
rlabel metal2 s 36174 79200 36230 80000 6 la_data_out[50]
port 396 nsew signal output
rlabel metal2 s 36450 79200 36506 80000 6 la_data_out[51]
port 397 nsew signal output
rlabel metal2 s 36726 79200 36782 80000 6 la_data_out[52]
port 398 nsew signal output
rlabel metal2 s 37002 79200 37058 80000 6 la_data_out[53]
port 399 nsew signal output
rlabel metal2 s 37278 79200 37334 80000 6 la_data_out[54]
port 400 nsew signal output
rlabel metal2 s 37554 79200 37610 80000 6 la_data_out[55]
port 401 nsew signal output
rlabel metal2 s 37830 79200 37886 80000 6 la_data_out[56]
port 402 nsew signal output
rlabel metal2 s 38106 79200 38162 80000 6 la_data_out[57]
port 403 nsew signal output
rlabel metal2 s 38382 79200 38438 80000 6 la_data_out[58]
port 404 nsew signal output
rlabel metal2 s 38658 79200 38714 80000 6 la_data_out[59]
port 405 nsew signal output
rlabel metal2 s 23754 79200 23810 80000 6 la_data_out[5]
port 406 nsew signal output
rlabel metal2 s 38934 79200 38990 80000 6 la_data_out[60]
port 407 nsew signal output
rlabel metal2 s 39210 79200 39266 80000 6 la_data_out[61]
port 408 nsew signal output
rlabel metal2 s 39486 79200 39542 80000 6 la_data_out[62]
port 409 nsew signal output
rlabel metal2 s 39762 79200 39818 80000 6 la_data_out[63]
port 410 nsew signal output
rlabel metal2 s 40038 79200 40094 80000 6 la_data_out[64]
port 411 nsew signal output
rlabel metal2 s 40314 79200 40370 80000 6 la_data_out[65]
port 412 nsew signal output
rlabel metal2 s 40590 79200 40646 80000 6 la_data_out[66]
port 413 nsew signal output
rlabel metal2 s 40866 79200 40922 80000 6 la_data_out[67]
port 414 nsew signal output
rlabel metal2 s 41142 79200 41198 80000 6 la_data_out[68]
port 415 nsew signal output
rlabel metal2 s 41418 79200 41474 80000 6 la_data_out[69]
port 416 nsew signal output
rlabel metal2 s 24030 79200 24086 80000 6 la_data_out[6]
port 417 nsew signal output
rlabel metal2 s 41694 79200 41750 80000 6 la_data_out[70]
port 418 nsew signal output
rlabel metal2 s 41970 79200 42026 80000 6 la_data_out[71]
port 419 nsew signal output
rlabel metal2 s 42246 79200 42302 80000 6 la_data_out[72]
port 420 nsew signal output
rlabel metal2 s 42522 79200 42578 80000 6 la_data_out[73]
port 421 nsew signal output
rlabel metal2 s 42798 79200 42854 80000 6 la_data_out[74]
port 422 nsew signal output
rlabel metal2 s 43074 79200 43130 80000 6 la_data_out[75]
port 423 nsew signal output
rlabel metal2 s 43350 79200 43406 80000 6 la_data_out[76]
port 424 nsew signal output
rlabel metal2 s 43626 79200 43682 80000 6 la_data_out[77]
port 425 nsew signal output
rlabel metal2 s 43902 79200 43958 80000 6 la_data_out[78]
port 426 nsew signal output
rlabel metal2 s 44178 79200 44234 80000 6 la_data_out[79]
port 427 nsew signal output
rlabel metal2 s 24306 79200 24362 80000 6 la_data_out[7]
port 428 nsew signal output
rlabel metal2 s 44454 79200 44510 80000 6 la_data_out[80]
port 429 nsew signal output
rlabel metal2 s 44730 79200 44786 80000 6 la_data_out[81]
port 430 nsew signal output
rlabel metal2 s 45006 79200 45062 80000 6 la_data_out[82]
port 431 nsew signal output
rlabel metal2 s 45282 79200 45338 80000 6 la_data_out[83]
port 432 nsew signal output
rlabel metal2 s 45558 79200 45614 80000 6 la_data_out[84]
port 433 nsew signal output
rlabel metal2 s 45834 79200 45890 80000 6 la_data_out[85]
port 434 nsew signal output
rlabel metal2 s 46110 79200 46166 80000 6 la_data_out[86]
port 435 nsew signal output
rlabel metal2 s 46386 79200 46442 80000 6 la_data_out[87]
port 436 nsew signal output
rlabel metal2 s 46662 79200 46718 80000 6 la_data_out[88]
port 437 nsew signal output
rlabel metal2 s 46938 79200 46994 80000 6 la_data_out[89]
port 438 nsew signal output
rlabel metal2 s 24582 79200 24638 80000 6 la_data_out[8]
port 439 nsew signal output
rlabel metal2 s 47214 79200 47270 80000 6 la_data_out[90]
port 440 nsew signal output
rlabel metal2 s 47490 79200 47546 80000 6 la_data_out[91]
port 441 nsew signal output
rlabel metal2 s 47766 79200 47822 80000 6 la_data_out[92]
port 442 nsew signal output
rlabel metal2 s 48042 79200 48098 80000 6 la_data_out[93]
port 443 nsew signal output
rlabel metal2 s 48318 79200 48374 80000 6 la_data_out[94]
port 444 nsew signal output
rlabel metal2 s 48594 79200 48650 80000 6 la_data_out[95]
port 445 nsew signal output
rlabel metal2 s 48870 79200 48926 80000 6 la_data_out[96]
port 446 nsew signal output
rlabel metal2 s 49146 79200 49202 80000 6 la_data_out[97]
port 447 nsew signal output
rlabel metal2 s 49422 79200 49478 80000 6 la_data_out[98]
port 448 nsew signal output
rlabel metal2 s 49698 79200 49754 80000 6 la_data_out[99]
port 449 nsew signal output
rlabel metal2 s 24858 79200 24914 80000 6 la_data_out[9]
port 450 nsew signal output
rlabel metal2 s 22466 79200 22522 80000 6 la_oenb[0]
port 451 nsew signal input
rlabel metal2 s 50066 79200 50122 80000 6 la_oenb[100]
port 452 nsew signal input
rlabel metal2 s 50342 79200 50398 80000 6 la_oenb[101]
port 453 nsew signal input
rlabel metal2 s 50618 79200 50674 80000 6 la_oenb[102]
port 454 nsew signal input
rlabel metal2 s 50894 79200 50950 80000 6 la_oenb[103]
port 455 nsew signal input
rlabel metal2 s 51170 79200 51226 80000 6 la_oenb[104]
port 456 nsew signal input
rlabel metal2 s 51446 79200 51502 80000 6 la_oenb[105]
port 457 nsew signal input
rlabel metal2 s 51722 79200 51778 80000 6 la_oenb[106]
port 458 nsew signal input
rlabel metal2 s 51998 79200 52054 80000 6 la_oenb[107]
port 459 nsew signal input
rlabel metal2 s 52274 79200 52330 80000 6 la_oenb[108]
port 460 nsew signal input
rlabel metal2 s 52550 79200 52606 80000 6 la_oenb[109]
port 461 nsew signal input
rlabel metal2 s 25226 79200 25282 80000 6 la_oenb[10]
port 462 nsew signal input
rlabel metal2 s 52826 79200 52882 80000 6 la_oenb[110]
port 463 nsew signal input
rlabel metal2 s 53102 79200 53158 80000 6 la_oenb[111]
port 464 nsew signal input
rlabel metal2 s 53378 79200 53434 80000 6 la_oenb[112]
port 465 nsew signal input
rlabel metal2 s 53654 79200 53710 80000 6 la_oenb[113]
port 466 nsew signal input
rlabel metal2 s 53930 79200 53986 80000 6 la_oenb[114]
port 467 nsew signal input
rlabel metal2 s 54206 79200 54262 80000 6 la_oenb[115]
port 468 nsew signal input
rlabel metal2 s 54482 79200 54538 80000 6 la_oenb[116]
port 469 nsew signal input
rlabel metal2 s 54758 79200 54814 80000 6 la_oenb[117]
port 470 nsew signal input
rlabel metal2 s 55034 79200 55090 80000 6 la_oenb[118]
port 471 nsew signal input
rlabel metal2 s 55310 79200 55366 80000 6 la_oenb[119]
port 472 nsew signal input
rlabel metal2 s 25502 79200 25558 80000 6 la_oenb[11]
port 473 nsew signal input
rlabel metal2 s 55586 79200 55642 80000 6 la_oenb[120]
port 474 nsew signal input
rlabel metal2 s 55862 79200 55918 80000 6 la_oenb[121]
port 475 nsew signal input
rlabel metal2 s 56138 79200 56194 80000 6 la_oenb[122]
port 476 nsew signal input
rlabel metal2 s 56414 79200 56470 80000 6 la_oenb[123]
port 477 nsew signal input
rlabel metal2 s 56690 79200 56746 80000 6 la_oenb[124]
port 478 nsew signal input
rlabel metal2 s 56966 79200 57022 80000 6 la_oenb[125]
port 479 nsew signal input
rlabel metal2 s 57242 79200 57298 80000 6 la_oenb[126]
port 480 nsew signal input
rlabel metal2 s 57518 79200 57574 80000 6 la_oenb[127]
port 481 nsew signal input
rlabel metal2 s 25778 79200 25834 80000 6 la_oenb[12]
port 482 nsew signal input
rlabel metal2 s 26054 79200 26110 80000 6 la_oenb[13]
port 483 nsew signal input
rlabel metal2 s 26330 79200 26386 80000 6 la_oenb[14]
port 484 nsew signal input
rlabel metal2 s 26606 79200 26662 80000 6 la_oenb[15]
port 485 nsew signal input
rlabel metal2 s 26882 79200 26938 80000 6 la_oenb[16]
port 486 nsew signal input
rlabel metal2 s 27158 79200 27214 80000 6 la_oenb[17]
port 487 nsew signal input
rlabel metal2 s 27434 79200 27490 80000 6 la_oenb[18]
port 488 nsew signal input
rlabel metal2 s 27710 79200 27766 80000 6 la_oenb[19]
port 489 nsew signal input
rlabel metal2 s 22742 79200 22798 80000 6 la_oenb[1]
port 490 nsew signal input
rlabel metal2 s 27986 79200 28042 80000 6 la_oenb[20]
port 491 nsew signal input
rlabel metal2 s 28262 79200 28318 80000 6 la_oenb[21]
port 492 nsew signal input
rlabel metal2 s 28538 79200 28594 80000 6 la_oenb[22]
port 493 nsew signal input
rlabel metal2 s 28814 79200 28870 80000 6 la_oenb[23]
port 494 nsew signal input
rlabel metal2 s 29090 79200 29146 80000 6 la_oenb[24]
port 495 nsew signal input
rlabel metal2 s 29366 79200 29422 80000 6 la_oenb[25]
port 496 nsew signal input
rlabel metal2 s 29642 79200 29698 80000 6 la_oenb[26]
port 497 nsew signal input
rlabel metal2 s 29918 79200 29974 80000 6 la_oenb[27]
port 498 nsew signal input
rlabel metal2 s 30194 79200 30250 80000 6 la_oenb[28]
port 499 nsew signal input
rlabel metal2 s 30470 79200 30526 80000 6 la_oenb[29]
port 500 nsew signal input
rlabel metal2 s 23018 79200 23074 80000 6 la_oenb[2]
port 501 nsew signal input
rlabel metal2 s 30746 79200 30802 80000 6 la_oenb[30]
port 502 nsew signal input
rlabel metal2 s 31022 79200 31078 80000 6 la_oenb[31]
port 503 nsew signal input
rlabel metal2 s 31298 79200 31354 80000 6 la_oenb[32]
port 504 nsew signal input
rlabel metal2 s 31574 79200 31630 80000 6 la_oenb[33]
port 505 nsew signal input
rlabel metal2 s 31850 79200 31906 80000 6 la_oenb[34]
port 506 nsew signal input
rlabel metal2 s 32126 79200 32182 80000 6 la_oenb[35]
port 507 nsew signal input
rlabel metal2 s 32402 79200 32458 80000 6 la_oenb[36]
port 508 nsew signal input
rlabel metal2 s 32678 79200 32734 80000 6 la_oenb[37]
port 509 nsew signal input
rlabel metal2 s 32954 79200 33010 80000 6 la_oenb[38]
port 510 nsew signal input
rlabel metal2 s 33230 79200 33286 80000 6 la_oenb[39]
port 511 nsew signal input
rlabel metal2 s 23294 79200 23350 80000 6 la_oenb[3]
port 512 nsew signal input
rlabel metal2 s 33506 79200 33562 80000 6 la_oenb[40]
port 513 nsew signal input
rlabel metal2 s 33782 79200 33838 80000 6 la_oenb[41]
port 514 nsew signal input
rlabel metal2 s 34058 79200 34114 80000 6 la_oenb[42]
port 515 nsew signal input
rlabel metal2 s 34334 79200 34390 80000 6 la_oenb[43]
port 516 nsew signal input
rlabel metal2 s 34610 79200 34666 80000 6 la_oenb[44]
port 517 nsew signal input
rlabel metal2 s 34886 79200 34942 80000 6 la_oenb[45]
port 518 nsew signal input
rlabel metal2 s 35162 79200 35218 80000 6 la_oenb[46]
port 519 nsew signal input
rlabel metal2 s 35438 79200 35494 80000 6 la_oenb[47]
port 520 nsew signal input
rlabel metal2 s 35714 79200 35770 80000 6 la_oenb[48]
port 521 nsew signal input
rlabel metal2 s 35990 79200 36046 80000 6 la_oenb[49]
port 522 nsew signal input
rlabel metal2 s 23570 79200 23626 80000 6 la_oenb[4]
port 523 nsew signal input
rlabel metal2 s 36266 79200 36322 80000 6 la_oenb[50]
port 524 nsew signal input
rlabel metal2 s 36542 79200 36598 80000 6 la_oenb[51]
port 525 nsew signal input
rlabel metal2 s 36818 79200 36874 80000 6 la_oenb[52]
port 526 nsew signal input
rlabel metal2 s 37094 79200 37150 80000 6 la_oenb[53]
port 527 nsew signal input
rlabel metal2 s 37370 79200 37426 80000 6 la_oenb[54]
port 528 nsew signal input
rlabel metal2 s 37646 79200 37702 80000 6 la_oenb[55]
port 529 nsew signal input
rlabel metal2 s 37922 79200 37978 80000 6 la_oenb[56]
port 530 nsew signal input
rlabel metal2 s 38198 79200 38254 80000 6 la_oenb[57]
port 531 nsew signal input
rlabel metal2 s 38474 79200 38530 80000 6 la_oenb[58]
port 532 nsew signal input
rlabel metal2 s 38750 79200 38806 80000 6 la_oenb[59]
port 533 nsew signal input
rlabel metal2 s 23846 79200 23902 80000 6 la_oenb[5]
port 534 nsew signal input
rlabel metal2 s 39026 79200 39082 80000 6 la_oenb[60]
port 535 nsew signal input
rlabel metal2 s 39302 79200 39358 80000 6 la_oenb[61]
port 536 nsew signal input
rlabel metal2 s 39578 79200 39634 80000 6 la_oenb[62]
port 537 nsew signal input
rlabel metal2 s 39854 79200 39910 80000 6 la_oenb[63]
port 538 nsew signal input
rlabel metal2 s 40130 79200 40186 80000 6 la_oenb[64]
port 539 nsew signal input
rlabel metal2 s 40406 79200 40462 80000 6 la_oenb[65]
port 540 nsew signal input
rlabel metal2 s 40682 79200 40738 80000 6 la_oenb[66]
port 541 nsew signal input
rlabel metal2 s 40958 79200 41014 80000 6 la_oenb[67]
port 542 nsew signal input
rlabel metal2 s 41234 79200 41290 80000 6 la_oenb[68]
port 543 nsew signal input
rlabel metal2 s 41510 79200 41566 80000 6 la_oenb[69]
port 544 nsew signal input
rlabel metal2 s 24122 79200 24178 80000 6 la_oenb[6]
port 545 nsew signal input
rlabel metal2 s 41786 79200 41842 80000 6 la_oenb[70]
port 546 nsew signal input
rlabel metal2 s 42062 79200 42118 80000 6 la_oenb[71]
port 547 nsew signal input
rlabel metal2 s 42338 79200 42394 80000 6 la_oenb[72]
port 548 nsew signal input
rlabel metal2 s 42614 79200 42670 80000 6 la_oenb[73]
port 549 nsew signal input
rlabel metal2 s 42890 79200 42946 80000 6 la_oenb[74]
port 550 nsew signal input
rlabel metal2 s 43166 79200 43222 80000 6 la_oenb[75]
port 551 nsew signal input
rlabel metal2 s 43442 79200 43498 80000 6 la_oenb[76]
port 552 nsew signal input
rlabel metal2 s 43718 79200 43774 80000 6 la_oenb[77]
port 553 nsew signal input
rlabel metal2 s 43994 79200 44050 80000 6 la_oenb[78]
port 554 nsew signal input
rlabel metal2 s 44270 79200 44326 80000 6 la_oenb[79]
port 555 nsew signal input
rlabel metal2 s 24398 79200 24454 80000 6 la_oenb[7]
port 556 nsew signal input
rlabel metal2 s 44546 79200 44602 80000 6 la_oenb[80]
port 557 nsew signal input
rlabel metal2 s 44822 79200 44878 80000 6 la_oenb[81]
port 558 nsew signal input
rlabel metal2 s 45098 79200 45154 80000 6 la_oenb[82]
port 559 nsew signal input
rlabel metal2 s 45374 79200 45430 80000 6 la_oenb[83]
port 560 nsew signal input
rlabel metal2 s 45650 79200 45706 80000 6 la_oenb[84]
port 561 nsew signal input
rlabel metal2 s 45926 79200 45982 80000 6 la_oenb[85]
port 562 nsew signal input
rlabel metal2 s 46202 79200 46258 80000 6 la_oenb[86]
port 563 nsew signal input
rlabel metal2 s 46478 79200 46534 80000 6 la_oenb[87]
port 564 nsew signal input
rlabel metal2 s 46754 79200 46810 80000 6 la_oenb[88]
port 565 nsew signal input
rlabel metal2 s 47030 79200 47086 80000 6 la_oenb[89]
port 566 nsew signal input
rlabel metal2 s 24674 79200 24730 80000 6 la_oenb[8]
port 567 nsew signal input
rlabel metal2 s 47306 79200 47362 80000 6 la_oenb[90]
port 568 nsew signal input
rlabel metal2 s 47582 79200 47638 80000 6 la_oenb[91]
port 569 nsew signal input
rlabel metal2 s 47858 79200 47914 80000 6 la_oenb[92]
port 570 nsew signal input
rlabel metal2 s 48134 79200 48190 80000 6 la_oenb[93]
port 571 nsew signal input
rlabel metal2 s 48410 79200 48466 80000 6 la_oenb[94]
port 572 nsew signal input
rlabel metal2 s 48686 79200 48742 80000 6 la_oenb[95]
port 573 nsew signal input
rlabel metal2 s 48962 79200 49018 80000 6 la_oenb[96]
port 574 nsew signal input
rlabel metal2 s 49238 79200 49294 80000 6 la_oenb[97]
port 575 nsew signal input
rlabel metal2 s 49514 79200 49570 80000 6 la_oenb[98]
port 576 nsew signal input
rlabel metal2 s 49790 79200 49846 80000 6 la_oenb[99]
port 577 nsew signal input
rlabel metal2 s 24950 79200 25006 80000 6 la_oenb[9]
port 578 nsew signal input
rlabel metal2 s 11794 79200 11850 80000 6 m_io_in[0]
port 579 nsew signal input
rlabel metal2 s 14554 79200 14610 80000 6 m_io_in[10]
port 580 nsew signal input
rlabel metal2 s 14830 79200 14886 80000 6 m_io_in[11]
port 581 nsew signal input
rlabel metal2 s 15106 79200 15162 80000 6 m_io_in[12]
port 582 nsew signal input
rlabel metal2 s 15382 79200 15438 80000 6 m_io_in[13]
port 583 nsew signal input
rlabel metal2 s 15658 79200 15714 80000 6 m_io_in[14]
port 584 nsew signal input
rlabel metal2 s 15934 79200 15990 80000 6 m_io_in[15]
port 585 nsew signal input
rlabel metal2 s 16210 79200 16266 80000 6 m_io_in[16]
port 586 nsew signal input
rlabel metal2 s 16486 79200 16542 80000 6 m_io_in[17]
port 587 nsew signal input
rlabel metal2 s 16762 79200 16818 80000 6 m_io_in[18]
port 588 nsew signal input
rlabel metal2 s 17038 79200 17094 80000 6 m_io_in[19]
port 589 nsew signal input
rlabel metal2 s 12070 79200 12126 80000 6 m_io_in[1]
port 590 nsew signal input
rlabel metal2 s 17314 79200 17370 80000 6 m_io_in[20]
port 591 nsew signal input
rlabel metal2 s 17590 79200 17646 80000 6 m_io_in[21]
port 592 nsew signal input
rlabel metal2 s 17866 79200 17922 80000 6 m_io_in[22]
port 593 nsew signal input
rlabel metal2 s 18142 79200 18198 80000 6 m_io_in[23]
port 594 nsew signal input
rlabel metal2 s 18418 79200 18474 80000 6 m_io_in[24]
port 595 nsew signal input
rlabel metal2 s 18694 79200 18750 80000 6 m_io_in[25]
port 596 nsew signal input
rlabel metal2 s 18970 79200 19026 80000 6 m_io_in[26]
port 597 nsew signal input
rlabel metal2 s 19246 79200 19302 80000 6 m_io_in[27]
port 598 nsew signal input
rlabel metal2 s 19522 79200 19578 80000 6 m_io_in[28]
port 599 nsew signal input
rlabel metal2 s 19798 79200 19854 80000 6 m_io_in[29]
port 600 nsew signal input
rlabel metal2 s 12346 79200 12402 80000 6 m_io_in[2]
port 601 nsew signal input
rlabel metal2 s 20074 79200 20130 80000 6 m_io_in[30]
port 602 nsew signal input
rlabel metal2 s 20350 79200 20406 80000 6 m_io_in[31]
port 603 nsew signal input
rlabel metal2 s 20626 79200 20682 80000 6 m_io_in[32]
port 604 nsew signal input
rlabel metal2 s 20902 79200 20958 80000 6 m_io_in[33]
port 605 nsew signal input
rlabel metal2 s 21178 79200 21234 80000 6 m_io_in[34]
port 606 nsew signal input
rlabel metal2 s 21454 79200 21510 80000 6 m_io_in[35]
port 607 nsew signal input
rlabel metal2 s 21730 79200 21786 80000 6 m_io_in[36]
port 608 nsew signal input
rlabel metal2 s 22006 79200 22062 80000 6 m_io_in[37]
port 609 nsew signal input
rlabel metal2 s 12622 79200 12678 80000 6 m_io_in[3]
port 610 nsew signal input
rlabel metal2 s 12898 79200 12954 80000 6 m_io_in[4]
port 611 nsew signal input
rlabel metal2 s 13174 79200 13230 80000 6 m_io_in[5]
port 612 nsew signal input
rlabel metal2 s 13450 79200 13506 80000 6 m_io_in[6]
port 613 nsew signal input
rlabel metal2 s 13726 79200 13782 80000 6 m_io_in[7]
port 614 nsew signal input
rlabel metal2 s 14002 79200 14058 80000 6 m_io_in[8]
port 615 nsew signal input
rlabel metal2 s 14278 79200 14334 80000 6 m_io_in[9]
port 616 nsew signal input
rlabel metal2 s 11886 79200 11942 80000 6 m_io_oeb[0]
port 617 nsew signal output
rlabel metal2 s 14646 79200 14702 80000 6 m_io_oeb[10]
port 618 nsew signal output
rlabel metal2 s 14922 79200 14978 80000 6 m_io_oeb[11]
port 619 nsew signal output
rlabel metal2 s 15198 79200 15254 80000 6 m_io_oeb[12]
port 620 nsew signal output
rlabel metal2 s 15474 79200 15530 80000 6 m_io_oeb[13]
port 621 nsew signal output
rlabel metal2 s 15750 79200 15806 80000 6 m_io_oeb[14]
port 622 nsew signal output
rlabel metal2 s 16026 79200 16082 80000 6 m_io_oeb[15]
port 623 nsew signal output
rlabel metal2 s 16302 79200 16358 80000 6 m_io_oeb[16]
port 624 nsew signal output
rlabel metal2 s 16578 79200 16634 80000 6 m_io_oeb[17]
port 625 nsew signal output
rlabel metal2 s 16854 79200 16910 80000 6 m_io_oeb[18]
port 626 nsew signal output
rlabel metal2 s 17130 79200 17186 80000 6 m_io_oeb[19]
port 627 nsew signal output
rlabel metal2 s 12162 79200 12218 80000 6 m_io_oeb[1]
port 628 nsew signal output
rlabel metal2 s 17406 79200 17462 80000 6 m_io_oeb[20]
port 629 nsew signal output
rlabel metal2 s 17682 79200 17738 80000 6 m_io_oeb[21]
port 630 nsew signal output
rlabel metal2 s 17958 79200 18014 80000 6 m_io_oeb[22]
port 631 nsew signal output
rlabel metal2 s 18234 79200 18290 80000 6 m_io_oeb[23]
port 632 nsew signal output
rlabel metal2 s 18510 79200 18566 80000 6 m_io_oeb[24]
port 633 nsew signal output
rlabel metal2 s 18786 79200 18842 80000 6 m_io_oeb[25]
port 634 nsew signal output
rlabel metal2 s 19062 79200 19118 80000 6 m_io_oeb[26]
port 635 nsew signal output
rlabel metal2 s 19338 79200 19394 80000 6 m_io_oeb[27]
port 636 nsew signal output
rlabel metal2 s 19614 79200 19670 80000 6 m_io_oeb[28]
port 637 nsew signal output
rlabel metal2 s 19890 79200 19946 80000 6 m_io_oeb[29]
port 638 nsew signal output
rlabel metal2 s 12438 79200 12494 80000 6 m_io_oeb[2]
port 639 nsew signal output
rlabel metal2 s 20166 79200 20222 80000 6 m_io_oeb[30]
port 640 nsew signal output
rlabel metal2 s 20442 79200 20498 80000 6 m_io_oeb[31]
port 641 nsew signal output
rlabel metal2 s 20718 79200 20774 80000 6 m_io_oeb[32]
port 642 nsew signal output
rlabel metal2 s 20994 79200 21050 80000 6 m_io_oeb[33]
port 643 nsew signal output
rlabel metal2 s 21270 79200 21326 80000 6 m_io_oeb[34]
port 644 nsew signal output
rlabel metal2 s 21546 79200 21602 80000 6 m_io_oeb[35]
port 645 nsew signal output
rlabel metal2 s 21822 79200 21878 80000 6 m_io_oeb[36]
port 646 nsew signal output
rlabel metal2 s 22098 79200 22154 80000 6 m_io_oeb[37]
port 647 nsew signal output
rlabel metal2 s 12714 79200 12770 80000 6 m_io_oeb[3]
port 648 nsew signal output
rlabel metal2 s 12990 79200 13046 80000 6 m_io_oeb[4]
port 649 nsew signal output
rlabel metal2 s 13266 79200 13322 80000 6 m_io_oeb[5]
port 650 nsew signal output
rlabel metal2 s 13542 79200 13598 80000 6 m_io_oeb[6]
port 651 nsew signal output
rlabel metal2 s 13818 79200 13874 80000 6 m_io_oeb[7]
port 652 nsew signal output
rlabel metal2 s 14094 79200 14150 80000 6 m_io_oeb[8]
port 653 nsew signal output
rlabel metal2 s 14370 79200 14426 80000 6 m_io_oeb[9]
port 654 nsew signal output
rlabel metal2 s 11978 79200 12034 80000 6 m_io_out[0]
port 655 nsew signal output
rlabel metal2 s 14738 79200 14794 80000 6 m_io_out[10]
port 656 nsew signal output
rlabel metal2 s 15014 79200 15070 80000 6 m_io_out[11]
port 657 nsew signal output
rlabel metal2 s 15290 79200 15346 80000 6 m_io_out[12]
port 658 nsew signal output
rlabel metal2 s 15566 79200 15622 80000 6 m_io_out[13]
port 659 nsew signal output
rlabel metal2 s 15842 79200 15898 80000 6 m_io_out[14]
port 660 nsew signal output
rlabel metal2 s 16118 79200 16174 80000 6 m_io_out[15]
port 661 nsew signal output
rlabel metal2 s 16394 79200 16450 80000 6 m_io_out[16]
port 662 nsew signal output
rlabel metal2 s 16670 79200 16726 80000 6 m_io_out[17]
port 663 nsew signal output
rlabel metal2 s 16946 79200 17002 80000 6 m_io_out[18]
port 664 nsew signal output
rlabel metal2 s 17222 79200 17278 80000 6 m_io_out[19]
port 665 nsew signal output
rlabel metal2 s 12254 79200 12310 80000 6 m_io_out[1]
port 666 nsew signal output
rlabel metal2 s 17498 79200 17554 80000 6 m_io_out[20]
port 667 nsew signal output
rlabel metal2 s 17774 79200 17830 80000 6 m_io_out[21]
port 668 nsew signal output
rlabel metal2 s 18050 79200 18106 80000 6 m_io_out[22]
port 669 nsew signal output
rlabel metal2 s 18326 79200 18382 80000 6 m_io_out[23]
port 670 nsew signal output
rlabel metal2 s 18602 79200 18658 80000 6 m_io_out[24]
port 671 nsew signal output
rlabel metal2 s 18878 79200 18934 80000 6 m_io_out[25]
port 672 nsew signal output
rlabel metal2 s 19154 79200 19210 80000 6 m_io_out[26]
port 673 nsew signal output
rlabel metal2 s 19430 79200 19486 80000 6 m_io_out[27]
port 674 nsew signal output
rlabel metal2 s 19706 79200 19762 80000 6 m_io_out[28]
port 675 nsew signal output
rlabel metal2 s 19982 79200 20038 80000 6 m_io_out[29]
port 676 nsew signal output
rlabel metal2 s 12530 79200 12586 80000 6 m_io_out[2]
port 677 nsew signal output
rlabel metal2 s 20258 79200 20314 80000 6 m_io_out[30]
port 678 nsew signal output
rlabel metal2 s 20534 79200 20590 80000 6 m_io_out[31]
port 679 nsew signal output
rlabel metal2 s 20810 79200 20866 80000 6 m_io_out[32]
port 680 nsew signal output
rlabel metal2 s 21086 79200 21142 80000 6 m_io_out[33]
port 681 nsew signal output
rlabel metal2 s 21362 79200 21418 80000 6 m_io_out[34]
port 682 nsew signal output
rlabel metal2 s 21638 79200 21694 80000 6 m_io_out[35]
port 683 nsew signal output
rlabel metal2 s 21914 79200 21970 80000 6 m_io_out[36]
port 684 nsew signal output
rlabel metal2 s 22190 79200 22246 80000 6 m_io_out[37]
port 685 nsew signal output
rlabel metal2 s 12806 79200 12862 80000 6 m_io_out[3]
port 686 nsew signal output
rlabel metal2 s 13082 79200 13138 80000 6 m_io_out[4]
port 687 nsew signal output
rlabel metal2 s 13358 79200 13414 80000 6 m_io_out[5]
port 688 nsew signal output
rlabel metal2 s 13634 79200 13690 80000 6 m_io_out[6]
port 689 nsew signal output
rlabel metal2 s 13910 79200 13966 80000 6 m_io_out[7]
port 690 nsew signal output
rlabel metal2 s 14186 79200 14242 80000 6 m_io_out[8]
port 691 nsew signal output
rlabel metal2 s 14462 79200 14518 80000 6 m_io_out[9]
port 692 nsew signal output
rlabel metal2 s 2042 79200 2098 80000 6 mgt_wb_ack_o
port 693 nsew signal output
rlabel metal2 s 2594 79200 2650 80000 6 mgt_wb_adr_i[0]
port 694 nsew signal input
rlabel metal2 s 5722 79200 5778 80000 6 mgt_wb_adr_i[10]
port 695 nsew signal input
rlabel metal2 s 5998 79200 6054 80000 6 mgt_wb_adr_i[11]
port 696 nsew signal input
rlabel metal2 s 6274 79200 6330 80000 6 mgt_wb_adr_i[12]
port 697 nsew signal input
rlabel metal2 s 6550 79200 6606 80000 6 mgt_wb_adr_i[13]
port 698 nsew signal input
rlabel metal2 s 6826 79200 6882 80000 6 mgt_wb_adr_i[14]
port 699 nsew signal input
rlabel metal2 s 7102 79200 7158 80000 6 mgt_wb_adr_i[15]
port 700 nsew signal input
rlabel metal2 s 7378 79200 7434 80000 6 mgt_wb_adr_i[16]
port 701 nsew signal input
rlabel metal2 s 7654 79200 7710 80000 6 mgt_wb_adr_i[17]
port 702 nsew signal input
rlabel metal2 s 7930 79200 7986 80000 6 mgt_wb_adr_i[18]
port 703 nsew signal input
rlabel metal2 s 8206 79200 8262 80000 6 mgt_wb_adr_i[19]
port 704 nsew signal input
rlabel metal2 s 2962 79200 3018 80000 6 mgt_wb_adr_i[1]
port 705 nsew signal input
rlabel metal2 s 8482 79200 8538 80000 6 mgt_wb_adr_i[20]
port 706 nsew signal input
rlabel metal2 s 8758 79200 8814 80000 6 mgt_wb_adr_i[21]
port 707 nsew signal input
rlabel metal2 s 9034 79200 9090 80000 6 mgt_wb_adr_i[22]
port 708 nsew signal input
rlabel metal2 s 9310 79200 9366 80000 6 mgt_wb_adr_i[23]
port 709 nsew signal input
rlabel metal2 s 9586 79200 9642 80000 6 mgt_wb_adr_i[24]
port 710 nsew signal input
rlabel metal2 s 9862 79200 9918 80000 6 mgt_wb_adr_i[25]
port 711 nsew signal input
rlabel metal2 s 10138 79200 10194 80000 6 mgt_wb_adr_i[26]
port 712 nsew signal input
rlabel metal2 s 10414 79200 10470 80000 6 mgt_wb_adr_i[27]
port 713 nsew signal input
rlabel metal2 s 10690 79200 10746 80000 6 mgt_wb_adr_i[28]
port 714 nsew signal input
rlabel metal2 s 10966 79200 11022 80000 6 mgt_wb_adr_i[29]
port 715 nsew signal input
rlabel metal2 s 3330 79200 3386 80000 6 mgt_wb_adr_i[2]
port 716 nsew signal input
rlabel metal2 s 11242 79200 11298 80000 6 mgt_wb_adr_i[30]
port 717 nsew signal input
rlabel metal2 s 11518 79200 11574 80000 6 mgt_wb_adr_i[31]
port 718 nsew signal input
rlabel metal2 s 3698 79200 3754 80000 6 mgt_wb_adr_i[3]
port 719 nsew signal input
rlabel metal2 s 4066 79200 4122 80000 6 mgt_wb_adr_i[4]
port 720 nsew signal input
rlabel metal2 s 4342 79200 4398 80000 6 mgt_wb_adr_i[5]
port 721 nsew signal input
rlabel metal2 s 4618 79200 4674 80000 6 mgt_wb_adr_i[6]
port 722 nsew signal input
rlabel metal2 s 4894 79200 4950 80000 6 mgt_wb_adr_i[7]
port 723 nsew signal input
rlabel metal2 s 5170 79200 5226 80000 6 mgt_wb_adr_i[8]
port 724 nsew signal input
rlabel metal2 s 5446 79200 5502 80000 6 mgt_wb_adr_i[9]
port 725 nsew signal input
rlabel metal2 s 2134 79200 2190 80000 6 mgt_wb_clk_i
port 726 nsew signal input
rlabel metal2 s 2226 79200 2282 80000 6 mgt_wb_cyc_i
port 727 nsew signal input
rlabel metal2 s 2686 79200 2742 80000 6 mgt_wb_dat_i[0]
port 728 nsew signal input
rlabel metal2 s 5814 79200 5870 80000 6 mgt_wb_dat_i[10]
port 729 nsew signal input
rlabel metal2 s 6090 79200 6146 80000 6 mgt_wb_dat_i[11]
port 730 nsew signal input
rlabel metal2 s 6366 79200 6422 80000 6 mgt_wb_dat_i[12]
port 731 nsew signal input
rlabel metal2 s 6642 79200 6698 80000 6 mgt_wb_dat_i[13]
port 732 nsew signal input
rlabel metal2 s 6918 79200 6974 80000 6 mgt_wb_dat_i[14]
port 733 nsew signal input
rlabel metal2 s 7194 79200 7250 80000 6 mgt_wb_dat_i[15]
port 734 nsew signal input
rlabel metal2 s 7470 79200 7526 80000 6 mgt_wb_dat_i[16]
port 735 nsew signal input
rlabel metal2 s 7746 79200 7802 80000 6 mgt_wb_dat_i[17]
port 736 nsew signal input
rlabel metal2 s 8022 79200 8078 80000 6 mgt_wb_dat_i[18]
port 737 nsew signal input
rlabel metal2 s 8298 79200 8354 80000 6 mgt_wb_dat_i[19]
port 738 nsew signal input
rlabel metal2 s 3054 79200 3110 80000 6 mgt_wb_dat_i[1]
port 739 nsew signal input
rlabel metal2 s 8574 79200 8630 80000 6 mgt_wb_dat_i[20]
port 740 nsew signal input
rlabel metal2 s 8850 79200 8906 80000 6 mgt_wb_dat_i[21]
port 741 nsew signal input
rlabel metal2 s 9126 79200 9182 80000 6 mgt_wb_dat_i[22]
port 742 nsew signal input
rlabel metal2 s 9402 79200 9458 80000 6 mgt_wb_dat_i[23]
port 743 nsew signal input
rlabel metal2 s 9678 79200 9734 80000 6 mgt_wb_dat_i[24]
port 744 nsew signal input
rlabel metal2 s 9954 79200 10010 80000 6 mgt_wb_dat_i[25]
port 745 nsew signal input
rlabel metal2 s 10230 79200 10286 80000 6 mgt_wb_dat_i[26]
port 746 nsew signal input
rlabel metal2 s 10506 79200 10562 80000 6 mgt_wb_dat_i[27]
port 747 nsew signal input
rlabel metal2 s 10782 79200 10838 80000 6 mgt_wb_dat_i[28]
port 748 nsew signal input
rlabel metal2 s 11058 79200 11114 80000 6 mgt_wb_dat_i[29]
port 749 nsew signal input
rlabel metal2 s 3422 79200 3478 80000 6 mgt_wb_dat_i[2]
port 750 nsew signal input
rlabel metal2 s 11334 79200 11390 80000 6 mgt_wb_dat_i[30]
port 751 nsew signal input
rlabel metal2 s 11610 79200 11666 80000 6 mgt_wb_dat_i[31]
port 752 nsew signal input
rlabel metal2 s 3790 79200 3846 80000 6 mgt_wb_dat_i[3]
port 753 nsew signal input
rlabel metal2 s 4158 79200 4214 80000 6 mgt_wb_dat_i[4]
port 754 nsew signal input
rlabel metal2 s 4434 79200 4490 80000 6 mgt_wb_dat_i[5]
port 755 nsew signal input
rlabel metal2 s 4710 79200 4766 80000 6 mgt_wb_dat_i[6]
port 756 nsew signal input
rlabel metal2 s 4986 79200 5042 80000 6 mgt_wb_dat_i[7]
port 757 nsew signal input
rlabel metal2 s 5262 79200 5318 80000 6 mgt_wb_dat_i[8]
port 758 nsew signal input
rlabel metal2 s 5538 79200 5594 80000 6 mgt_wb_dat_i[9]
port 759 nsew signal input
rlabel metal2 s 2778 79200 2834 80000 6 mgt_wb_dat_o[0]
port 760 nsew signal output
rlabel metal2 s 5906 79200 5962 80000 6 mgt_wb_dat_o[10]
port 761 nsew signal output
rlabel metal2 s 6182 79200 6238 80000 6 mgt_wb_dat_o[11]
port 762 nsew signal output
rlabel metal2 s 6458 79200 6514 80000 6 mgt_wb_dat_o[12]
port 763 nsew signal output
rlabel metal2 s 6734 79200 6790 80000 6 mgt_wb_dat_o[13]
port 764 nsew signal output
rlabel metal2 s 7010 79200 7066 80000 6 mgt_wb_dat_o[14]
port 765 nsew signal output
rlabel metal2 s 7286 79200 7342 80000 6 mgt_wb_dat_o[15]
port 766 nsew signal output
rlabel metal2 s 7562 79200 7618 80000 6 mgt_wb_dat_o[16]
port 767 nsew signal output
rlabel metal2 s 7838 79200 7894 80000 6 mgt_wb_dat_o[17]
port 768 nsew signal output
rlabel metal2 s 8114 79200 8170 80000 6 mgt_wb_dat_o[18]
port 769 nsew signal output
rlabel metal2 s 8390 79200 8446 80000 6 mgt_wb_dat_o[19]
port 770 nsew signal output
rlabel metal2 s 3146 79200 3202 80000 6 mgt_wb_dat_o[1]
port 771 nsew signal output
rlabel metal2 s 8666 79200 8722 80000 6 mgt_wb_dat_o[20]
port 772 nsew signal output
rlabel metal2 s 8942 79200 8998 80000 6 mgt_wb_dat_o[21]
port 773 nsew signal output
rlabel metal2 s 9218 79200 9274 80000 6 mgt_wb_dat_o[22]
port 774 nsew signal output
rlabel metal2 s 9494 79200 9550 80000 6 mgt_wb_dat_o[23]
port 775 nsew signal output
rlabel metal2 s 9770 79200 9826 80000 6 mgt_wb_dat_o[24]
port 776 nsew signal output
rlabel metal2 s 10046 79200 10102 80000 6 mgt_wb_dat_o[25]
port 777 nsew signal output
rlabel metal2 s 10322 79200 10378 80000 6 mgt_wb_dat_o[26]
port 778 nsew signal output
rlabel metal2 s 10598 79200 10654 80000 6 mgt_wb_dat_o[27]
port 779 nsew signal output
rlabel metal2 s 10874 79200 10930 80000 6 mgt_wb_dat_o[28]
port 780 nsew signal output
rlabel metal2 s 11150 79200 11206 80000 6 mgt_wb_dat_o[29]
port 781 nsew signal output
rlabel metal2 s 3514 79200 3570 80000 6 mgt_wb_dat_o[2]
port 782 nsew signal output
rlabel metal2 s 11426 79200 11482 80000 6 mgt_wb_dat_o[30]
port 783 nsew signal output
rlabel metal2 s 11702 79200 11758 80000 6 mgt_wb_dat_o[31]
port 784 nsew signal output
rlabel metal2 s 3882 79200 3938 80000 6 mgt_wb_dat_o[3]
port 785 nsew signal output
rlabel metal2 s 4250 79200 4306 80000 6 mgt_wb_dat_o[4]
port 786 nsew signal output
rlabel metal2 s 4526 79200 4582 80000 6 mgt_wb_dat_o[5]
port 787 nsew signal output
rlabel metal2 s 4802 79200 4858 80000 6 mgt_wb_dat_o[6]
port 788 nsew signal output
rlabel metal2 s 5078 79200 5134 80000 6 mgt_wb_dat_o[7]
port 789 nsew signal output
rlabel metal2 s 5354 79200 5410 80000 6 mgt_wb_dat_o[8]
port 790 nsew signal output
rlabel metal2 s 5630 79200 5686 80000 6 mgt_wb_dat_o[9]
port 791 nsew signal output
rlabel metal2 s 2318 79200 2374 80000 6 mgt_wb_rst_i
port 792 nsew signal input
rlabel metal2 s 2870 79200 2926 80000 6 mgt_wb_sel_i[0]
port 793 nsew signal input
rlabel metal2 s 3238 79200 3294 80000 6 mgt_wb_sel_i[1]
port 794 nsew signal input
rlabel metal2 s 3606 79200 3662 80000 6 mgt_wb_sel_i[2]
port 795 nsew signal input
rlabel metal2 s 3974 79200 4030 80000 6 mgt_wb_sel_i[3]
port 796 nsew signal input
rlabel metal2 s 2410 79200 2466 80000 6 mgt_wb_stb_i
port 797 nsew signal input
rlabel metal2 s 2502 79200 2558 80000 6 mgt_wb_we_i
port 798 nsew signal input
rlabel metal2 s 57886 79200 57942 80000 6 user_clock2
port 799 nsew signal input
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 800 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 800 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 801 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 801 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8374198
string GDS_FILE /home/piotro/caravel_user_project/openlane/interconnect_outer/runs/22_12_30_12_19/results/signoff/interconnect_outer.magic.gds
string GDS_START 760442
<< end >>

